-- q_sys.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity q_sys is
	port (
		clock_bridge_0_in_clk_clk               : in    std_logic                    := '0';             --               clock_bridge_0_in_clk.clk
		enet_clk_125m_in_clk                    : in    std_logic                    := '0';             --                    enet_clk_125m_in.clk
		enet_pll_areset_conduit_export          : in    std_logic                    := '0';             --             enet_pll_areset_conduit.export
		enet_pll_c0_125m_clk                    : out   std_logic;                                       --                    enet_pll_c0_125m.clk
		enet_pll_c1_25m_clk                     : out   std_logic;                                       --                     enet_pll_c1_25m.clk
		enet_pll_c2_2m5_clk                     : out   std_logic;                                       --                     enet_pll_c2_2m5.clk
		enet_pll_c3_125m_shift_clk              : out   std_logic;                                       --              enet_pll_c3_125m_shift.clk
		enet_pll_c4_25m_shift_clk               : out   std_logic;                                       --               enet_pll_c4_25m_shift.clk
		enet_pll_locked_conduit_export          : out   std_logic;                                       --             enet_pll_locked_conduit.export
		eth_tse_mac_mdio_connection_mdc         : out   std_logic;                                       --         eth_tse_mac_mdio_connection.mdc
		eth_tse_mac_mdio_connection_mdio_in     : in    std_logic                    := '0';             --                                    .mdio_in
		eth_tse_mac_mdio_connection_mdio_out    : out   std_logic;                                       --                                    .mdio_out
		eth_tse_mac_mdio_connection_mdio_oen    : out   std_logic;                                       --                                    .mdio_oen
		eth_tse_mac_rgmii_connection_rgmii_in   : in    std_logic_vector(3 downto 0) := (others => '0'); --        eth_tse_mac_rgmii_connection.rgmii_in
		eth_tse_mac_rgmii_connection_rgmii_out  : out   std_logic_vector(3 downto 0);                    --                                    .rgmii_out
		eth_tse_mac_rgmii_connection_rx_control : in    std_logic                    := '0';             --                                    .rx_control
		eth_tse_mac_rgmii_connection_tx_control : out   std_logic;                                       --                                    .tx_control
		eth_tse_mac_status_connection_set_10    : in    std_logic                    := '0';             --       eth_tse_mac_status_connection.set_10
		eth_tse_mac_status_connection_set_1000  : in    std_logic                    := '0';             --                                    .set_1000
		eth_tse_mac_status_connection_eth_mode  : out   std_logic;                                       --                                    .eth_mode
		eth_tse_mac_status_connection_ena_10    : out   std_logic;                                       --                                    .ena_10
		eth_tse_pcs_mac_rx_clock_connection_clk : in    std_logic                    := '0';             -- eth_tse_pcs_mac_rx_clock_connection.clk
		eth_tse_pcs_mac_tx_clock_connection_clk : in    std_logic                    := '0';             -- eth_tse_pcs_mac_tx_clock_connection.clk
		hbus_clk_clk                            : in    std_logic                    := '0';             --                            hbus_clk.clk
		hbus_reset_reset_n                      : in    std_logic                    := '0';             --                          hbus_reset.reset_n
		hyperbus_controller_top_HB_RSTn         : out   std_logic;                                       --             hyperbus_controller_top.HB_RSTn
		hyperbus_controller_top_HB_CLK0         : out   std_logic;                                       --                                    .HB_CLK0
		hyperbus_controller_top_HB_CLK0n        : out   std_logic;                                       --                                    .HB_CLK0n
		hyperbus_controller_top_HB_CLK1         : out   std_logic;                                       --                                    .HB_CLK1
		hyperbus_controller_top_HB_CLK1n        : out   std_logic;                                       --                                    .HB_CLK1n
		hyperbus_controller_top_HB_CS0n         : out   std_logic;                                       --                                    .HB_CS0n
		hyperbus_controller_top_HB_CS1n         : out   std_logic;                                       --                                    .HB_CS1n
		hyperbus_controller_top_HB_WPn          : out   std_logic;                                       --                                    .HB_WPn
		hyperbus_controller_top_HB_RWDS         : inout std_logic                    := '0';             --                                    .HB_RWDS
		hyperbus_controller_top_HB_dq           : inout std_logic_vector(7 downto 0) := (others => '0'); --                                    .HB_dq
		hyperbus_controller_top_HB_RSTOn        : in    std_logic                    := '0';             --                                    .HB_RSTOn
		hyperbus_controller_top_HB_INTn         : in    std_logic                    := '0';             --                                    .HB_INTn
		led_pio_external_connection_export      : out   std_logic_vector(3 downto 0);                    --         led_pio_external_connection.export
		opencores_i2c_scl_pad_io                : inout std_logic                    := '0';             --                       opencores_i2c.scl_pad_io
		opencores_i2c_sda_pad_io                : inout std_logic                    := '0';             --                                    .sda_pad_io
		reset_enet_reset_n                      : in    std_logic                    := '0';             --                          reset_enet.reset_n
		user_dipsw_external_connection_export   : in    std_logic_vector(3 downto 0) := (others => '0'); --      user_dipsw_external_connection.export
		user_pb_external_connection_export      : in    std_logic_vector(3 downto 0) := (others => '0')  --         user_pb_external_connection.export
	);
end entity q_sys;

architecture rtl of q_sys is
	component q_sys_cpu is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(26 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_burstcount                        : out std_logic_vector(3 downto 0);                     -- burstcount
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(26 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_burstcount                        : out std_logic_vector(3 downto 0);                     -- burstcount
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component q_sys_cpu;

	component q_sys_descriptor_memory is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(10 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component q_sys_descriptor_memory;

	component q_sys_enet_pll is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			read               : in  std_logic                     := 'X';             -- read
			write              : in  std_logic                     := 'X';             -- write
			address            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0                 : out std_logic;                                        -- clk
			c1                 : out std_logic;                                        -- clk
			c2                 : out std_logic;                                        -- clk
			c3                 : out std_logic;                                        -- clk
			c4                 : out std_logic;                                        -- clk
			areset             : in  std_logic                     := 'X';             -- export
			locked             : out std_logic;                                        -- export
			scandone           : out std_logic;                                        -- export
			scandataout        : out std_logic;                                        -- export
			phasedone          : out std_logic;                                        -- export
			phasecounterselect : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			phaseupdown        : in  std_logic                     := 'X';             -- export
			phasestep          : in  std_logic                     := 'X';             -- export
			scanclk            : in  std_logic                     := 'X';             -- export
			scanclkena         : in  std_logic                     := 'X';             -- export
			scandata           : in  std_logic                     := 'X';             -- export
			configupdate       : in  std_logic                     := 'X'              -- export
		);
	end component q_sys_enet_pll;

	component q_sys_eth_tse is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset         : in  std_logic                     := 'X';             -- reset
			reg_addr      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			reg_data_out  : out std_logic_vector(31 downto 0);                    -- readdata
			reg_rd        : in  std_logic                     := 'X';             -- read
			reg_data_in   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			reg_wr        : in  std_logic                     := 'X';             -- write
			reg_busy      : out std_logic;                                        -- waitrequest
			tx_clk        : in  std_logic                     := 'X';             -- clk
			rx_clk        : in  std_logic                     := 'X';             -- clk
			set_10        : in  std_logic                     := 'X';             -- set_10
			set_1000      : in  std_logic                     := 'X';             -- set_1000
			eth_mode      : out std_logic;                                        -- eth_mode
			ena_10        : out std_logic;                                        -- ena_10
			rgmii_in      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- rgmii_in
			rgmii_out     : out std_logic_vector(3 downto 0);                     -- rgmii_out
			rx_control    : in  std_logic                     := 'X';             -- rx_control
			tx_control    : out std_logic;                                        -- tx_control
			ff_rx_clk     : in  std_logic                     := 'X';             -- clk
			ff_tx_clk     : in  std_logic                     := 'X';             -- clk
			ff_rx_data    : out std_logic_vector(31 downto 0);                    -- data
			ff_rx_eop     : out std_logic;                                        -- endofpacket
			rx_err        : out std_logic_vector(5 downto 0);                     -- error
			ff_rx_mod     : out std_logic_vector(1 downto 0);                     -- empty
			ff_rx_rdy     : in  std_logic                     := 'X';             -- ready
			ff_rx_sop     : out std_logic;                                        -- startofpacket
			ff_rx_dval    : out std_logic;                                        -- valid
			ff_tx_data    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			ff_tx_eop     : in  std_logic                     := 'X';             -- endofpacket
			ff_tx_err     : in  std_logic                     := 'X';             -- error
			ff_tx_mod     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- empty
			ff_tx_rdy     : out std_logic;                                        -- ready
			ff_tx_sop     : in  std_logic                     := 'X';             -- startofpacket
			ff_tx_wren    : in  std_logic                     := 'X';             -- valid
			mdc           : out std_logic;                                        -- mdc
			mdio_in       : in  std_logic                     := 'X';             -- mdio_in
			mdio_out      : out std_logic;                                        -- mdio_out
			mdio_oen      : out std_logic;                                        -- mdio_oen
			magic_wakeup  : out std_logic;                                        -- magic_wakeup
			magic_sleep_n : in  std_logic                     := 'X';             -- magic_sleep_n
			ff_tx_crc_fwd : in  std_logic                     := 'X';             -- ff_tx_crc_fwd
			ff_tx_septy   : out std_logic;                                        -- ff_tx_septy
			tx_ff_uflow   : out std_logic;                                        -- tx_ff_uflow
			ff_tx_a_full  : out std_logic;                                        -- ff_tx_a_full
			ff_tx_a_empty : out std_logic;                                        -- ff_tx_a_empty
			rx_err_stat   : out std_logic_vector(17 downto 0);                    -- rx_err_stat
			rx_frm_type   : out std_logic_vector(3 downto 0);                     -- rx_frm_type
			ff_rx_dsav    : out std_logic;                                        -- ff_rx_dsav
			ff_rx_a_full  : out std_logic;                                        -- ff_rx_a_full
			ff_rx_a_empty : out std_logic                                         -- ff_rx_a_empty
		);
	end component q_sys_eth_tse;

	component q_sys_ext_epcq_flash is
		generic (
			DEVICE_FAMILY     : string  := "";
			ASI_WIDTH         : integer := 1;
			CS_WIDTH          : integer := 1;
			ADDR_WIDTH        : integer := 19;
			ASMI_ADDR_WIDTH   : integer := 24;
			ENABLE_4BYTE_ADDR : integer := 0;
			CHIP_SELS         : integer := 1
		);
		port (
			avl_csr_read         : in  std_logic                     := 'X';             -- read
			avl_csr_waitrequest  : out std_logic;                                        -- waitrequest
			avl_csr_write        : in  std_logic                     := 'X';             -- write
			avl_csr_addr         : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			avl_csr_wrdata       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avl_csr_rddata       : out std_logic_vector(31 downto 0);                    -- readdata
			avl_csr_rddata_valid : out std_logic;                                        -- readdatavalid
			avl_mem_write        : in  std_logic                     := 'X';             -- write
			avl_mem_burstcount   : in  std_logic_vector(6 downto 0)  := (others => 'X'); -- burstcount
			avl_mem_waitrequest  : out std_logic;                                        -- waitrequest
			avl_mem_read         : in  std_logic                     := 'X';             -- read
			avl_mem_addr         : in  std_logic_vector(20 downto 0) := (others => 'X'); -- address
			avl_mem_wrdata       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avl_mem_rddata       : out std_logic_vector(31 downto 0);                    -- readdata
			avl_mem_rddata_valid : out std_logic;                                        -- readdatavalid
			avl_mem_byteenable   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			irq                  : out std_logic;                                        -- irq
			clk                  : in  std_logic                     := 'X';             -- clk
			reset_n              : in  std_logic                     := 'X'              -- reset_n
		);
	end component q_sys_ext_epcq_flash;

	component q_sys_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component q_sys_jtag_uart;

	component q_sys_led_pio is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(3 downto 0)                      -- export
		);
	end component q_sys_led_pio;

	component altera_avalon_mm_bridge is
		generic (
			DATA_WIDTH        : integer := 32;
			SYMBOL_WIDTH      : integer := 8;
			HDL_ADDR_WIDTH    : integer := 10;
			BURSTCOUNT_WIDTH  : integer := 1;
			PIPELINE_COMMAND  : integer := 1;
			PIPELINE_RESPONSE : integer := 1
		);
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			reset            : in  std_logic                     := 'X';             -- reset
			s0_waitrequest   : out std_logic;                                        -- waitrequest
			s0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                        -- readdatavalid
			s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			s0_address       : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			s0_write         : in  std_logic                     := 'X';             -- write
			s0_read          : in  std_logic                     := 'X';             -- read
			s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			s0_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			m0_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			m0_burstcount    : out std_logic_vector(0 downto 0);                     -- burstcount
			m0_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			m0_address       : out std_logic_vector(14 downto 0);                    -- address
			m0_write         : out std_logic;                                        -- write
			m0_read          : out std_logic;                                        -- read
			m0_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess   : out std_logic;                                        -- debugaccess
			s0_response      : out std_logic_vector(1 downto 0);                     -- response
			m0_response      : in  std_logic_vector(1 downto 0)  := (others => 'X')  -- response
		);
	end component altera_avalon_mm_bridge;

	component q_sys_msgdma_rx is
		port (
			mm_write_address                           : out std_logic_vector(26 downto 0);                    -- address
			mm_write_write                             : out std_logic;                                        -- write
			mm_write_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			mm_write_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			mm_write_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			descriptor_read_master_address             : out std_logic_vector(14 downto 0);                    -- address
			descriptor_read_master_read                : out std_logic;                                        -- read
			descriptor_read_master_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			descriptor_read_master_waitrequest         : in  std_logic                     := 'X';             -- waitrequest
			descriptor_read_master_readdatavalid       : in  std_logic                     := 'X';             -- readdatavalid
			descriptor_write_master_address            : out std_logic_vector(14 downto 0);                    -- address
			descriptor_write_master_write              : out std_logic;                                        -- write
			descriptor_write_master_byteenable         : out std_logic_vector(3 downto 0);                     -- byteenable
			descriptor_write_master_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			descriptor_write_master_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			descriptor_write_master_response           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			descriptor_write_master_writeresponsevalid : in  std_logic                     := 'X';             -- writeresponsevalid
			clock_clk                                  : in  std_logic                     := 'X';             -- clk
			reset_n_reset_n                            : in  std_logic                     := 'X';             -- reset_n
			csr_writedata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			csr_write                                  : in  std_logic                     := 'X';             -- write
			csr_byteenable                             : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			csr_readdata                               : out std_logic_vector(31 downto 0);                    -- readdata
			csr_read                                   : in  std_logic                     := 'X';             -- read
			csr_address                                : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			prefetcher_csr_address                     : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			prefetcher_csr_read                        : in  std_logic                     := 'X';             -- read
			prefetcher_csr_write                       : in  std_logic                     := 'X';             -- write
			prefetcher_csr_writedata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			prefetcher_csr_readdata                    : out std_logic_vector(31 downto 0);                    -- readdata
			csr_irq_irq                                : out std_logic;                                        -- irq
			st_sink_data                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			st_sink_valid                              : in  std_logic                     := 'X';             -- valid
			st_sink_ready                              : out std_logic;                                        -- ready
			st_sink_startofpacket                      : in  std_logic                     := 'X';             -- startofpacket
			st_sink_endofpacket                        : in  std_logic                     := 'X';             -- endofpacket
			st_sink_empty                              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- empty
			st_sink_error                              : in  std_logic_vector(5 downto 0)  := (others => 'X')  -- error
		);
	end component q_sys_msgdma_rx;

	component q_sys_msgdma_tx is
		port (
			mm_read_address                            : out std_logic_vector(26 downto 0);                    -- address
			mm_read_read                               : out std_logic;                                        -- read
			mm_read_byteenable                         : out std_logic_vector(3 downto 0);                     -- byteenable
			mm_read_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			mm_read_waitrequest                        : in  std_logic                     := 'X';             -- waitrequest
			mm_read_readdatavalid                      : in  std_logic                     := 'X';             -- readdatavalid
			descriptor_read_master_address             : out std_logic_vector(14 downto 0);                    -- address
			descriptor_read_master_read                : out std_logic;                                        -- read
			descriptor_read_master_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			descriptor_read_master_waitrequest         : in  std_logic                     := 'X';             -- waitrequest
			descriptor_read_master_readdatavalid       : in  std_logic                     := 'X';             -- readdatavalid
			descriptor_write_master_address            : out std_logic_vector(14 downto 0);                    -- address
			descriptor_write_master_write              : out std_logic;                                        -- write
			descriptor_write_master_byteenable         : out std_logic_vector(3 downto 0);                     -- byteenable
			descriptor_write_master_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			descriptor_write_master_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			descriptor_write_master_response           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			descriptor_write_master_writeresponsevalid : in  std_logic                     := 'X';             -- writeresponsevalid
			clock_clk                                  : in  std_logic                     := 'X';             -- clk
			reset_n_reset_n                            : in  std_logic                     := 'X';             -- reset_n
			csr_writedata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			csr_write                                  : in  std_logic                     := 'X';             -- write
			csr_byteenable                             : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			csr_readdata                               : out std_logic_vector(31 downto 0);                    -- readdata
			csr_read                                   : in  std_logic                     := 'X';             -- read
			csr_address                                : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			prefetcher_csr_address                     : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			prefetcher_csr_read                        : in  std_logic                     := 'X';             -- read
			prefetcher_csr_write                       : in  std_logic                     := 'X';             -- write
			prefetcher_csr_writedata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			prefetcher_csr_readdata                    : out std_logic_vector(31 downto 0);                    -- readdata
			csr_irq_irq                                : out std_logic;                                        -- irq
			st_source_data                             : out std_logic_vector(31 downto 0);                    -- data
			st_source_valid                            : out std_logic;                                        -- valid
			st_source_ready                            : in  std_logic                     := 'X';             -- ready
			st_source_startofpacket                    : out std_logic;                                        -- startofpacket
			st_source_endofpacket                      : out std_logic;                                        -- endofpacket
			st_source_empty                            : out std_logic_vector(1 downto 0);                     -- empty
			st_source_error                            : out std_logic                                         -- error
		);
	end component q_sys_msgdma_tx;

	component q_sys_onchip_ram is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component q_sys_onchip_ram;

	component opencores_i2c is
		generic (
			FIXED_PRESCALE : integer := 0
		);
		port (
			wb_clk_i   : in    std_logic                    := 'X';             -- clk
			wb_rst_i   : in    std_logic                    := 'X';             -- reset
			scl_pad_io : inout std_logic                    := 'X';             -- export
			sda_pad_io : inout std_logic                    := 'X';             -- export
			wb_adr_i   : in    std_logic_vector(2 downto 0) := (others => 'X'); -- address
			wb_dat_i   : in    std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			wb_dat_o   : out   std_logic_vector(7 downto 0);                    -- readdata
			wb_we_i    : in    std_logic                    := 'X';             -- write
			wb_stb_i   : in    std_logic                    := 'X';             -- chipselect
			wb_ack_o   : out   std_logic;                                       -- waitrequest_n
			wb_inta_o  : out   std_logic                                        -- irq
		);
	end component opencores_i2c;

	component q_sys_remote_update is
		port (
			avl_csr_write         : in  std_logic                     := 'X';             -- write
			avl_csr_read          : in  std_logic                     := 'X';             -- read
			avl_csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avl_csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			avl_csr_readdatavalid : out std_logic;                                        -- readdatavalid
			avl_csr_waitrequest   : out std_logic;                                        -- waitrequest
			avl_csr_address       : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- address
			clock_clk             : in  std_logic                     := 'X';             -- clk
			reset_reset           : in  std_logic                     := 'X'              -- reset
		);
	end component q_sys_remote_update;

	component sll_hyperbus_controller_top is
		generic (
			g_iavs0_addr_width         : integer                       := 18;
			g_iavs0_data_width         : integer                       := 32;
			g_iavs0_av_numsymbols      : integer                       := 4;
			g_iavs0_burstcount_width   : integer                       := 1;
			g_iavs0_linewrap_burst     : integer                       := 0;
			g_iavs0_register_rdata     : integer                       := 0;
			g_iavs0_register_wdata     : integer                       := 0;
			g_include_reg_avalon       : integer                       := 0;
			g_include_internal_pll     : integer                       := 1;
			g_input_clk_freq_in_mhz    : integer                       := 0;
			g_hyperbus_freq_in_mhz     : integer                       := 0;
			g_iavs_freq_in_mhz         : integer                       := 0;
			g_same_iavs_hyperbus_clk   : integer                       := 0;
			g_config_rd_buffer_as_sram : integer                       := 1;
			g_config_wr_buffer_as_sram : integer                       := 1;
			g_device_family            : string                        := "MAX 10";
			g_num_chipselect           : integer                       := 0;
			g_dev0_config              : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			g_dev1_config              : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			g_dev0_timing              : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			g_dev1_timing              : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			g_include_dual_rwds_pin    : integer                       := 0;
			g_dqin_rdata_width         : integer                       := 8
		);
		port (
			in_clk               : in    std_logic                     := 'X';             -- clk
			i_ext_rstn           : in    std_logic                     := 'X';             -- reset_n
			i_iavs0_clk          : in    std_logic                     := 'X';             -- clk
			i_iavs0_rstn         : in    std_logic                     := 'X';             -- reset_n
			i_iavs0_addr         : in    std_logic_vector(21 downto 0) := (others => 'X'); -- address
			i_iavs0_burstcount   : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- burstcount
			o_iavs0_wait_request : out   std_logic;                                        -- waitrequest
			i_iavs0_do_wr        : in    std_logic                     := 'X';             -- write
			i_iavs0_byteenable   : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			i_iavs0_wdata        : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			i_iavs0_do_rd        : in    std_logic                     := 'X';             -- read
			o_iavs0_rdata        : out   std_logic_vector(31 downto 0);                    -- readdata
			o_iavs0_rdata_valid  : out   std_logic;                                        -- readdatavalid
			HB_RSTn              : out   std_logic;                                        -- HB_RSTn
			HB_CLK0              : out   std_logic;                                        -- HB_CLK0
			HB_CLK0n             : out   std_logic;                                        -- HB_CLK0n
			HB_CLK1              : out   std_logic;                                        -- HB_CLK1
			HB_CLK1n             : out   std_logic;                                        -- HB_CLK1n
			HB_CS0n              : out   std_logic;                                        -- HB_CS0n
			HB_CS1n              : out   std_logic;                                        -- HB_CS1n
			HB_WPn               : out   std_logic;                                        -- HB_WPn
			HB_RWDS              : inout std_logic                     := 'X';             -- HB_RWDS
			HB_dq                : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- HB_dq
			HB_RSTOn             : in    std_logic                     := 'X';             -- HB_RSTOn
			HB_INTn              : in    std_logic                     := 'X';             -- HB_INTn
			o_av_out_clk         : out   std_logic;                                        -- clk
			o_av_out_rstn        : out   std_logic;                                        -- reset_n
			o_iavs0_resp         : out   std_logic_vector(1 downto 0);                     -- response
			i_iavsr_addr         : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			i_iavsr_do_wr        : in    std_logic                     := 'X';             -- write
			i_iavsr_do_rd        : in    std_logic                     := 'X';             -- read
			i_iavsr_wdata        : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			o_iavsr_rdata        : out   std_logic_vector(31 downto 0)                     -- readdata
		);
	end component sll_hyperbus_controller_top;

	component q_sys_sys_clk_timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component q_sys_sys_clk_timer;

	component q_sys_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component q_sys_sysid;

	component q_sys_user_dipsw is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(3 downto 0)  := (others => 'X')  -- export
		);
	end component q_sys_user_dipsw;

	component userhw is
		port (
			clk       : in  std_logic                     := 'X';             -- clk
			read      : in  std_logic                     := 'X';             -- read
			write     : in  std_logic                     := 'X';             -- write
			address   : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata  : out std_logic_vector(31 downto 0);                    -- readdata
			rst       : in  std_logic                     := 'X'              -- reset
		);
	end component userhw;

	component q_sys_mm_interconnect_0 is
		port (
			clock_bridge_0_out_clk_clk                                             : in  std_logic                     := 'X';             -- clk
			sll_hyperbus_controller_top_0_o_av_out_clk_clk                         : in  std_logic                     := 'X';             -- clk
			cpu_reset_reset_bridge_in_reset_reset                                  : in  std_logic                     := 'X';             -- reset
			ext_epcq_flash_reset_reset_bridge_in_reset_reset                       : in  std_logic                     := 'X';             -- reset
			sll_hyperbus_controller_top_0_i_iavs0_rstn_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			cpu_data_master_address                                                : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			cpu_data_master_waitrequest                                            : out std_logic;                                        -- waitrequest
			cpu_data_master_burstcount                                             : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- burstcount
			cpu_data_master_byteenable                                             : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_data_master_read                                                   : in  std_logic                     := 'X';             -- read
			cpu_data_master_readdata                                               : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_data_master_readdatavalid                                          : out std_logic;                                        -- readdatavalid
			cpu_data_master_write                                                  : in  std_logic                     := 'X';             -- write
			cpu_data_master_writedata                                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_data_master_debugaccess                                            : in  std_logic                     := 'X';             -- debugaccess
			cpu_instruction_master_address                                         : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			cpu_instruction_master_waitrequest                                     : out std_logic;                                        -- waitrequest
			cpu_instruction_master_burstcount                                      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- burstcount
			cpu_instruction_master_read                                            : in  std_logic                     := 'X';             -- read
			cpu_instruction_master_readdata                                        : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_instruction_master_readdatavalid                                   : out std_logic;                                        -- readdatavalid
			msgdma_rx_mm_write_address                                             : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			msgdma_rx_mm_write_waitrequest                                         : out std_logic;                                        -- waitrequest
			msgdma_rx_mm_write_byteenable                                          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			msgdma_rx_mm_write_write                                               : in  std_logic                     := 'X';             -- write
			msgdma_rx_mm_write_writedata                                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			msgdma_tx_mm_read_address                                              : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			msgdma_tx_mm_read_waitrequest                                          : out std_logic;                                        -- waitrequest
			msgdma_tx_mm_read_byteenable                                           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			msgdma_tx_mm_read_read                                                 : in  std_logic                     := 'X';             -- read
			msgdma_tx_mm_read_readdata                                             : out std_logic_vector(31 downto 0);                    -- readdata
			msgdma_tx_mm_read_readdatavalid                                        : out std_logic;                                        -- readdatavalid
			cpu_debug_mem_slave_address                                            : out std_logic_vector(8 downto 0);                     -- address
			cpu_debug_mem_slave_write                                              : out std_logic;                                        -- write
			cpu_debug_mem_slave_read                                               : out std_logic;                                        -- read
			cpu_debug_mem_slave_readdata                                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_debug_mem_slave_writedata                                          : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_debug_mem_slave_byteenable                                         : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_debug_mem_slave_waitrequest                                        : in  std_logic                     := 'X';             -- waitrequest
			cpu_debug_mem_slave_debugaccess                                        : out std_logic;                                        -- debugaccess
			ext_epcq_flash_avl_csr_address                                         : out std_logic_vector(3 downto 0);                     -- address
			ext_epcq_flash_avl_csr_write                                           : out std_logic;                                        -- write
			ext_epcq_flash_avl_csr_read                                            : out std_logic;                                        -- read
			ext_epcq_flash_avl_csr_readdata                                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ext_epcq_flash_avl_csr_writedata                                       : out std_logic_vector(31 downto 0);                    -- writedata
			ext_epcq_flash_avl_csr_readdatavalid                                   : in  std_logic                     := 'X';             -- readdatavalid
			ext_epcq_flash_avl_csr_waitrequest                                     : in  std_logic                     := 'X';             -- waitrequest
			ext_epcq_flash_avl_mem_address                                         : out std_logic_vector(20 downto 0);                    -- address
			ext_epcq_flash_avl_mem_write                                           : out std_logic;                                        -- write
			ext_epcq_flash_avl_mem_read                                            : out std_logic;                                        -- read
			ext_epcq_flash_avl_mem_readdata                                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ext_epcq_flash_avl_mem_writedata                                       : out std_logic_vector(31 downto 0);                    -- writedata
			ext_epcq_flash_avl_mem_burstcount                                      : out std_logic_vector(6 downto 0);                     -- burstcount
			ext_epcq_flash_avl_mem_byteenable                                      : out std_logic_vector(3 downto 0);                     -- byteenable
			ext_epcq_flash_avl_mem_readdatavalid                                   : in  std_logic                     := 'X';             -- readdatavalid
			ext_epcq_flash_avl_mem_waitrequest                                     : in  std_logic                     := 'X';             -- waitrequest
			mm_bridge_0_s0_address                                                 : out std_logic_vector(14 downto 0);                    -- address
			mm_bridge_0_s0_write                                                   : out std_logic;                                        -- write
			mm_bridge_0_s0_read                                                    : out std_logic;                                        -- read
			mm_bridge_0_s0_readdata                                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			mm_bridge_0_s0_writedata                                               : out std_logic_vector(31 downto 0);                    -- writedata
			mm_bridge_0_s0_burstcount                                              : out std_logic_vector(0 downto 0);                     -- burstcount
			mm_bridge_0_s0_byteenable                                              : out std_logic_vector(3 downto 0);                     -- byteenable
			mm_bridge_0_s0_readdatavalid                                           : in  std_logic                     := 'X';             -- readdatavalid
			mm_bridge_0_s0_waitrequest                                             : in  std_logic                     := 'X';             -- waitrequest
			mm_bridge_0_s0_debugaccess                                             : out std_logic;                                        -- debugaccess
			onchip_ram_s1_address                                                  : out std_logic_vector(8 downto 0);                     -- address
			onchip_ram_s1_write                                                    : out std_logic;                                        -- write
			onchip_ram_s1_readdata                                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_ram_s1_writedata                                                : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_ram_s1_byteenable                                               : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_ram_s1_chipselect                                               : out std_logic;                                        -- chipselect
			onchip_ram_s1_clken                                                    : out std_logic;                                        -- clken
			remote_update_avl_csr_address                                          : out std_logic_vector(4 downto 0);                     -- address
			remote_update_avl_csr_write                                            : out std_logic;                                        -- write
			remote_update_avl_csr_read                                             : out std_logic;                                        -- read
			remote_update_avl_csr_readdata                                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			remote_update_avl_csr_writedata                                        : out std_logic_vector(31 downto 0);                    -- writedata
			remote_update_avl_csr_readdatavalid                                    : in  std_logic                     := 'X';             -- readdatavalid
			remote_update_avl_csr_waitrequest                                      : in  std_logic                     := 'X';             -- waitrequest
			sll_hyperbus_controller_top_0_iavs0_address                            : out std_logic_vector(21 downto 0);                    -- address
			sll_hyperbus_controller_top_0_iavs0_write                              : out std_logic;                                        -- write
			sll_hyperbus_controller_top_0_iavs0_read                               : out std_logic;                                        -- read
			sll_hyperbus_controller_top_0_iavs0_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sll_hyperbus_controller_top_0_iavs0_writedata                          : out std_logic_vector(31 downto 0);                    -- writedata
			sll_hyperbus_controller_top_0_iavs0_burstcount                         : out std_logic_vector(3 downto 0);                     -- burstcount
			sll_hyperbus_controller_top_0_iavs0_byteenable                         : out std_logic_vector(3 downto 0);                     -- byteenable
			sll_hyperbus_controller_top_0_iavs0_readdatavalid                      : in  std_logic                     := 'X';             -- readdatavalid
			sll_hyperbus_controller_top_0_iavs0_waitrequest                        : in  std_logic                     := 'X'              -- waitrequest
		);
	end component q_sys_mm_interconnect_0;

	component q_sys_mm_interconnect_1 is
		port (
			sll_hyperbus_controller_top_0_o_av_out_clk_clk       : in  std_logic                     := 'X';             -- clk
			descriptor_memory_reset1_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			msgdma_rx_reset_n_reset_bridge_in_reset_reset        : in  std_logic                     := 'X';             -- reset
			mm_bridge_0_m0_address                               : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			mm_bridge_0_m0_waitrequest                           : out std_logic;                                        -- waitrequest
			mm_bridge_0_m0_burstcount                            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			mm_bridge_0_m0_byteenable                            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			mm_bridge_0_m0_read                                  : in  std_logic                     := 'X';             -- read
			mm_bridge_0_m0_readdata                              : out std_logic_vector(31 downto 0);                    -- readdata
			mm_bridge_0_m0_readdatavalid                         : out std_logic;                                        -- readdatavalid
			mm_bridge_0_m0_write                                 : in  std_logic                     := 'X';             -- write
			mm_bridge_0_m0_writedata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			mm_bridge_0_m0_debugaccess                           : in  std_logic                     := 'X';             -- debugaccess
			msgdma_rx_descriptor_read_master_address             : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			msgdma_rx_descriptor_read_master_waitrequest         : out std_logic;                                        -- waitrequest
			msgdma_rx_descriptor_read_master_read                : in  std_logic                     := 'X';             -- read
			msgdma_rx_descriptor_read_master_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			msgdma_rx_descriptor_read_master_readdatavalid       : out std_logic;                                        -- readdatavalid
			msgdma_rx_descriptor_write_master_address            : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			msgdma_rx_descriptor_write_master_waitrequest        : out std_logic;                                        -- waitrequest
			msgdma_rx_descriptor_write_master_byteenable         : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			msgdma_rx_descriptor_write_master_write              : in  std_logic                     := 'X';             -- write
			msgdma_rx_descriptor_write_master_writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			msgdma_rx_descriptor_write_master_response           : out std_logic_vector(1 downto 0);                     -- response
			msgdma_rx_descriptor_write_master_writeresponsevalid : out std_logic;                                        -- writeresponsevalid
			msgdma_tx_descriptor_read_master_address             : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			msgdma_tx_descriptor_read_master_waitrequest         : out std_logic;                                        -- waitrequest
			msgdma_tx_descriptor_read_master_read                : in  std_logic                     := 'X';             -- read
			msgdma_tx_descriptor_read_master_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			msgdma_tx_descriptor_read_master_readdatavalid       : out std_logic;                                        -- readdatavalid
			msgdma_tx_descriptor_write_master_address            : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			msgdma_tx_descriptor_write_master_waitrequest        : out std_logic;                                        -- waitrequest
			msgdma_tx_descriptor_write_master_byteenable         : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			msgdma_tx_descriptor_write_master_write              : in  std_logic                     := 'X';             -- write
			msgdma_tx_descriptor_write_master_writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			msgdma_tx_descriptor_write_master_response           : out std_logic_vector(1 downto 0);                     -- response
			msgdma_tx_descriptor_write_master_writeresponsevalid : out std_logic;                                        -- writeresponsevalid
			descriptor_memory_s1_address                         : out std_logic_vector(10 downto 0);                    -- address
			descriptor_memory_s1_write                           : out std_logic;                                        -- write
			descriptor_memory_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			descriptor_memory_s1_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			descriptor_memory_s1_byteenable                      : out std_logic_vector(3 downto 0);                     -- byteenable
			descriptor_memory_s1_chipselect                      : out std_logic;                                        -- chipselect
			descriptor_memory_s1_clken                           : out std_logic;                                        -- clken
			eth_tse_control_port_address                         : out std_logic_vector(7 downto 0);                     -- address
			eth_tse_control_port_write                           : out std_logic;                                        -- write
			eth_tse_control_port_read                            : out std_logic;                                        -- read
			eth_tse_control_port_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			eth_tse_control_port_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			eth_tse_control_port_waitrequest                     : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_address                  : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write                    : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read                     : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata                : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest              : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect               : out std_logic;                                        -- chipselect
			led_pio_s1_address                                   : out std_logic_vector(1 downto 0);                     -- address
			led_pio_s1_write                                     : out std_logic;                                        -- write
			led_pio_s1_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			led_pio_s1_writedata                                 : out std_logic_vector(31 downto 0);                    -- writedata
			led_pio_s1_chipselect                                : out std_logic;                                        -- chipselect
			msgdma_rx_csr_address                                : out std_logic_vector(2 downto 0);                     -- address
			msgdma_rx_csr_write                                  : out std_logic;                                        -- write
			msgdma_rx_csr_read                                   : out std_logic;                                        -- read
			msgdma_rx_csr_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			msgdma_rx_csr_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			msgdma_rx_csr_byteenable                             : out std_logic_vector(3 downto 0);                     -- byteenable
			msgdma_rx_prefetcher_csr_address                     : out std_logic_vector(2 downto 0);                     -- address
			msgdma_rx_prefetcher_csr_write                       : out std_logic;                                        -- write
			msgdma_rx_prefetcher_csr_read                        : out std_logic;                                        -- read
			msgdma_rx_prefetcher_csr_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			msgdma_rx_prefetcher_csr_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			msgdma_tx_csr_address                                : out std_logic_vector(2 downto 0);                     -- address
			msgdma_tx_csr_write                                  : out std_logic;                                        -- write
			msgdma_tx_csr_read                                   : out std_logic;                                        -- read
			msgdma_tx_csr_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			msgdma_tx_csr_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			msgdma_tx_csr_byteenable                             : out std_logic_vector(3 downto 0);                     -- byteenable
			msgdma_tx_prefetcher_csr_address                     : out std_logic_vector(2 downto 0);                     -- address
			msgdma_tx_prefetcher_csr_write                       : out std_logic;                                        -- write
			msgdma_tx_prefetcher_csr_read                        : out std_logic;                                        -- read
			msgdma_tx_prefetcher_csr_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			msgdma_tx_prefetcher_csr_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			opencores_i2c_0_avalon_slave_0_address               : out std_logic_vector(2 downto 0);                     -- address
			opencores_i2c_0_avalon_slave_0_write                 : out std_logic;                                        -- write
			opencores_i2c_0_avalon_slave_0_readdata              : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			opencores_i2c_0_avalon_slave_0_writedata             : out std_logic_vector(7 downto 0);                     -- writedata
			opencores_i2c_0_avalon_slave_0_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			opencores_i2c_0_avalon_slave_0_chipselect            : out std_logic;                                        -- chipselect
			sys_clk_timer_s1_address                             : out std_logic_vector(2 downto 0);                     -- address
			sys_clk_timer_s1_write                               : out std_logic;                                        -- write
			sys_clk_timer_s1_readdata                            : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sys_clk_timer_s1_writedata                           : out std_logic_vector(15 downto 0);                    -- writedata
			sys_clk_timer_s1_chipselect                          : out std_logic;                                        -- chipselect
			sysid_control_slave_address                          : out std_logic_vector(0 downto 0);                     -- address
			sysid_control_slave_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			user_dipsw_s1_address                                : out std_logic_vector(1 downto 0);                     -- address
			user_dipsw_s1_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			user_pb_s1_address                                   : out std_logic_vector(1 downto 0);                     -- address
			user_pb_s1_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			userhw_0_avalon_slave_0_address                      : out std_logic_vector(2 downto 0);                     -- address
			userhw_0_avalon_slave_0_write                        : out std_logic;                                        -- write
			userhw_0_avalon_slave_0_read                         : out std_logic;                                        -- read
			userhw_0_avalon_slave_0_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			userhw_0_avalon_slave_0_writedata                    : out std_logic_vector(31 downto 0)                     -- writedata
		);
	end component q_sys_mm_interconnect_1;

	component q_sys_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component q_sys_irq_mapper;

	component q_sys_avalon_st_adapter is
		generic (
			inBitsPerSymbol : integer := 8;
			inUsePackets    : integer := 0;
			inDataWidth     : integer := 8;
			inChannelWidth  : integer := 3;
			inErrorWidth    : integer := 2;
			inUseEmptyPort  : integer := 0;
			inUseValid      : integer := 1;
			inUseReady      : integer := 1;
			inReadyLatency  : integer := 0;
			outDataWidth    : integer := 32;
			outChannelWidth : integer := 3;
			outErrorWidth   : integer := 2;
			outUseEmptyPort : integer := 0;
			outUseValid     : integer := 1;
			outUseReady     : integer := 1;
			outReadyLatency : integer := 0
		);
		port (
			in_clk_0_clk        : in  std_logic                     := 'X';             -- clk
			in_rst_0_reset      : in  std_logic                     := 'X';             -- reset
			in_0_data           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			in_0_valid          : in  std_logic                     := 'X';             -- valid
			in_0_ready          : out std_logic;                                        -- ready
			in_0_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_0_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			in_0_empty          : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- empty
			in_0_error          : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- error
			out_0_data          : out std_logic_vector(31 downto 0);                    -- data
			out_0_valid         : out std_logic;                                        -- valid
			out_0_ready         : in  std_logic                     := 'X';             -- ready
			out_0_startofpacket : out std_logic;                                        -- startofpacket
			out_0_endofpacket   : out std_logic;                                        -- endofpacket
			out_0_empty         : out std_logic_vector(1 downto 0);                     -- empty
			out_0_error         : out std_logic_vector(5 downto 0)                      -- error
		);
	end component q_sys_avalon_st_adapter;

	component q_sys_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component q_sys_rst_controller;

	component q_sys_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component q_sys_rst_controller_001;

	signal msgdma_tx_st_source_valid                                           : std_logic;                     -- msgdma_tx:st_source_valid -> eth_tse:ff_tx_wren
	signal msgdma_tx_st_source_data                                            : std_logic_vector(31 downto 0); -- msgdma_tx:st_source_data -> eth_tse:ff_tx_data
	signal msgdma_tx_st_source_ready                                           : std_logic;                     -- eth_tse:ff_tx_rdy -> msgdma_tx:st_source_ready
	signal msgdma_tx_st_source_startofpacket                                   : std_logic;                     -- msgdma_tx:st_source_startofpacket -> eth_tse:ff_tx_sop
	signal msgdma_tx_st_source_endofpacket                                     : std_logic;                     -- msgdma_tx:st_source_endofpacket -> eth_tse:ff_tx_eop
	signal msgdma_tx_st_source_error                                           : std_logic;                     -- msgdma_tx:st_source_error -> eth_tse:ff_tx_err
	signal msgdma_tx_st_source_empty                                           : std_logic_vector(1 downto 0);  -- msgdma_tx:st_source_empty -> eth_tse:ff_tx_mod
	signal sll_hyperbus_controller_top_0_o_av_out_clk_clk                      : std_logic;                     -- sll_hyperbus_controller_top_0:o_av_out_clk -> [avalon_st_adapter:in_clk_0_clk, cpu:clk, descriptor_memory:clk, eth_tse:clk, eth_tse:ff_rx_clk, eth_tse:ff_tx_clk, irq_mapper:clk, jtag_uart:clk, led_pio:clk, mm_bridge_0:clk, mm_interconnect_0:sll_hyperbus_controller_top_0_o_av_out_clk_clk, mm_interconnect_1:sll_hyperbus_controller_top_0_o_av_out_clk_clk, msgdma_rx:clock_clk, msgdma_tx:clock_clk, onchip_ram:clk, opencores_i2c_0:wb_clk_i, rst_controller:clk, sll_hyperbus_controller_top_0:i_iavs0_clk, sys_clk_timer:clk, sysid:clock, user_dipsw:clk, user_pb:clk, userhw_0:clk]
	signal sll_hyperbus_controller_top_0_o_av_out_rstn_reset                   : std_logic;                     -- sll_hyperbus_controller_top_0:o_av_out_rstn -> [msgdma_rx:reset_n_reset_n, msgdma_tx:reset_n_reset_n, sll_hyperbus_controller_top_0:i_iavs0_rstn, sll_hyperbus_controller_top_0_o_av_out_rstn_reset:in, user_dipsw:reset_n, user_pb:reset_n]
	signal cpu_data_master_readdata                                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	signal cpu_data_master_waitrequest                                         : std_logic;                     -- mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	signal cpu_data_master_debugaccess                                         : std_logic;                     -- cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	signal cpu_data_master_address                                             : std_logic_vector(26 downto 0); -- cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	signal cpu_data_master_byteenable                                          : std_logic_vector(3 downto 0);  -- cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	signal cpu_data_master_read                                                : std_logic;                     -- cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	signal cpu_data_master_readdatavalid                                       : std_logic;                     -- mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	signal cpu_data_master_write                                               : std_logic;                     -- cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	signal cpu_data_master_writedata                                           : std_logic_vector(31 downto 0); -- cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	signal cpu_data_master_burstcount                                          : std_logic_vector(3 downto 0);  -- cpu:d_burstcount -> mm_interconnect_0:cpu_data_master_burstcount
	signal cpu_instruction_master_readdata                                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	signal cpu_instruction_master_waitrequest                                  : std_logic;                     -- mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	signal cpu_instruction_master_address                                      : std_logic_vector(26 downto 0); -- cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	signal cpu_instruction_master_read                                         : std_logic;                     -- cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	signal cpu_instruction_master_readdatavalid                                : std_logic;                     -- mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	signal cpu_instruction_master_burstcount                                   : std_logic_vector(3 downto 0);  -- cpu:i_burstcount -> mm_interconnect_0:cpu_instruction_master_burstcount
	signal msgdma_tx_mm_read_readdata                                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:msgdma_tx_mm_read_readdata -> msgdma_tx:mm_read_readdata
	signal msgdma_tx_mm_read_waitrequest                                       : std_logic;                     -- mm_interconnect_0:msgdma_tx_mm_read_waitrequest -> msgdma_tx:mm_read_waitrequest
	signal msgdma_tx_mm_read_address                                           : std_logic_vector(26 downto 0); -- msgdma_tx:mm_read_address -> mm_interconnect_0:msgdma_tx_mm_read_address
	signal msgdma_tx_mm_read_read                                              : std_logic;                     -- msgdma_tx:mm_read_read -> mm_interconnect_0:msgdma_tx_mm_read_read
	signal msgdma_tx_mm_read_byteenable                                        : std_logic_vector(3 downto 0);  -- msgdma_tx:mm_read_byteenable -> mm_interconnect_0:msgdma_tx_mm_read_byteenable
	signal msgdma_tx_mm_read_readdatavalid                                     : std_logic;                     -- mm_interconnect_0:msgdma_tx_mm_read_readdatavalid -> msgdma_tx:mm_read_readdatavalid
	signal msgdma_rx_mm_write_waitrequest                                      : std_logic;                     -- mm_interconnect_0:msgdma_rx_mm_write_waitrequest -> msgdma_rx:mm_write_waitrequest
	signal msgdma_rx_mm_write_address                                          : std_logic_vector(26 downto 0); -- msgdma_rx:mm_write_address -> mm_interconnect_0:msgdma_rx_mm_write_address
	signal msgdma_rx_mm_write_byteenable                                       : std_logic_vector(3 downto 0);  -- msgdma_rx:mm_write_byteenable -> mm_interconnect_0:msgdma_rx_mm_write_byteenable
	signal msgdma_rx_mm_write_write                                            : std_logic;                     -- msgdma_rx:mm_write_write -> mm_interconnect_0:msgdma_rx_mm_write_write
	signal msgdma_rx_mm_write_writedata                                        : std_logic_vector(31 downto 0); -- msgdma_rx:mm_write_writedata -> mm_interconnect_0:msgdma_rx_mm_write_writedata
	signal mm_interconnect_0_ext_epcq_flash_avl_csr_readdata                   : std_logic_vector(31 downto 0); -- ext_epcq_flash:avl_csr_rddata -> mm_interconnect_0:ext_epcq_flash_avl_csr_readdata
	signal mm_interconnect_0_ext_epcq_flash_avl_csr_waitrequest                : std_logic;                     -- ext_epcq_flash:avl_csr_waitrequest -> mm_interconnect_0:ext_epcq_flash_avl_csr_waitrequest
	signal mm_interconnect_0_ext_epcq_flash_avl_csr_address                    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:ext_epcq_flash_avl_csr_address -> ext_epcq_flash:avl_csr_addr
	signal mm_interconnect_0_ext_epcq_flash_avl_csr_read                       : std_logic;                     -- mm_interconnect_0:ext_epcq_flash_avl_csr_read -> ext_epcq_flash:avl_csr_read
	signal mm_interconnect_0_ext_epcq_flash_avl_csr_readdatavalid              : std_logic;                     -- ext_epcq_flash:avl_csr_rddata_valid -> mm_interconnect_0:ext_epcq_flash_avl_csr_readdatavalid
	signal mm_interconnect_0_ext_epcq_flash_avl_csr_write                      : std_logic;                     -- mm_interconnect_0:ext_epcq_flash_avl_csr_write -> ext_epcq_flash:avl_csr_write
	signal mm_interconnect_0_ext_epcq_flash_avl_csr_writedata                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:ext_epcq_flash_avl_csr_writedata -> ext_epcq_flash:avl_csr_wrdata
	signal mm_interconnect_0_remote_update_avl_csr_readdata                    : std_logic_vector(31 downto 0); -- remote_update:avl_csr_readdata -> mm_interconnect_0:remote_update_avl_csr_readdata
	signal mm_interconnect_0_remote_update_avl_csr_waitrequest                 : std_logic;                     -- remote_update:avl_csr_waitrequest -> mm_interconnect_0:remote_update_avl_csr_waitrequest
	signal mm_interconnect_0_remote_update_avl_csr_address                     : std_logic_vector(4 downto 0);  -- mm_interconnect_0:remote_update_avl_csr_address -> remote_update:avl_csr_address
	signal mm_interconnect_0_remote_update_avl_csr_read                        : std_logic;                     -- mm_interconnect_0:remote_update_avl_csr_read -> remote_update:avl_csr_read
	signal mm_interconnect_0_remote_update_avl_csr_readdatavalid               : std_logic;                     -- remote_update:avl_csr_readdatavalid -> mm_interconnect_0:remote_update_avl_csr_readdatavalid
	signal mm_interconnect_0_remote_update_avl_csr_write                       : std_logic;                     -- mm_interconnect_0:remote_update_avl_csr_write -> remote_update:avl_csr_write
	signal mm_interconnect_0_remote_update_avl_csr_writedata                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:remote_update_avl_csr_writedata -> remote_update:avl_csr_writedata
	signal mm_interconnect_0_ext_epcq_flash_avl_mem_readdata                   : std_logic_vector(31 downto 0); -- ext_epcq_flash:avl_mem_rddata -> mm_interconnect_0:ext_epcq_flash_avl_mem_readdata
	signal mm_interconnect_0_ext_epcq_flash_avl_mem_waitrequest                : std_logic;                     -- ext_epcq_flash:avl_mem_waitrequest -> mm_interconnect_0:ext_epcq_flash_avl_mem_waitrequest
	signal mm_interconnect_0_ext_epcq_flash_avl_mem_address                    : std_logic_vector(20 downto 0); -- mm_interconnect_0:ext_epcq_flash_avl_mem_address -> ext_epcq_flash:avl_mem_addr
	signal mm_interconnect_0_ext_epcq_flash_avl_mem_read                       : std_logic;                     -- mm_interconnect_0:ext_epcq_flash_avl_mem_read -> ext_epcq_flash:avl_mem_read
	signal mm_interconnect_0_ext_epcq_flash_avl_mem_byteenable                 : std_logic_vector(3 downto 0);  -- mm_interconnect_0:ext_epcq_flash_avl_mem_byteenable -> ext_epcq_flash:avl_mem_byteenable
	signal mm_interconnect_0_ext_epcq_flash_avl_mem_readdatavalid              : std_logic;                     -- ext_epcq_flash:avl_mem_rddata_valid -> mm_interconnect_0:ext_epcq_flash_avl_mem_readdatavalid
	signal mm_interconnect_0_ext_epcq_flash_avl_mem_write                      : std_logic;                     -- mm_interconnect_0:ext_epcq_flash_avl_mem_write -> ext_epcq_flash:avl_mem_write
	signal mm_interconnect_0_ext_epcq_flash_avl_mem_writedata                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:ext_epcq_flash_avl_mem_writedata -> ext_epcq_flash:avl_mem_wrdata
	signal mm_interconnect_0_ext_epcq_flash_avl_mem_burstcount                 : std_logic_vector(6 downto 0);  -- mm_interconnect_0:ext_epcq_flash_avl_mem_burstcount -> ext_epcq_flash:avl_mem_burstcount
	signal mm_interconnect_0_cpu_debug_mem_slave_readdata                      : std_logic_vector(31 downto 0); -- cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_debug_mem_slave_waitrequest                   : std_logic;                     -- cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_debug_mem_slave_debugaccess                   : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_debug_mem_slave_address                       : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	signal mm_interconnect_0_cpu_debug_mem_slave_read                          : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	signal mm_interconnect_0_cpu_debug_mem_slave_byteenable                    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_debug_mem_slave_write                         : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	signal mm_interconnect_0_cpu_debug_mem_slave_writedata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	signal mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_readdata      : std_logic_vector(31 downto 0); -- sll_hyperbus_controller_top_0:o_iavs0_rdata -> mm_interconnect_0:sll_hyperbus_controller_top_0_iavs0_readdata
	signal mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_waitrequest   : std_logic;                     -- sll_hyperbus_controller_top_0:o_iavs0_wait_request -> mm_interconnect_0:sll_hyperbus_controller_top_0_iavs0_waitrequest
	signal mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_address       : std_logic_vector(21 downto 0); -- mm_interconnect_0:sll_hyperbus_controller_top_0_iavs0_address -> sll_hyperbus_controller_top_0:i_iavs0_addr
	signal mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_read          : std_logic;                     -- mm_interconnect_0:sll_hyperbus_controller_top_0_iavs0_read -> sll_hyperbus_controller_top_0:i_iavs0_do_rd
	signal mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_byteenable    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:sll_hyperbus_controller_top_0_iavs0_byteenable -> sll_hyperbus_controller_top_0:i_iavs0_byteenable
	signal mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_readdatavalid : std_logic;                     -- sll_hyperbus_controller_top_0:o_iavs0_rdata_valid -> mm_interconnect_0:sll_hyperbus_controller_top_0_iavs0_readdatavalid
	signal mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_write         : std_logic;                     -- mm_interconnect_0:sll_hyperbus_controller_top_0_iavs0_write -> sll_hyperbus_controller_top_0:i_iavs0_do_wr
	signal mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_writedata     : std_logic_vector(31 downto 0); -- mm_interconnect_0:sll_hyperbus_controller_top_0_iavs0_writedata -> sll_hyperbus_controller_top_0:i_iavs0_wdata
	signal mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_burstcount    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:sll_hyperbus_controller_top_0_iavs0_burstcount -> sll_hyperbus_controller_top_0:i_iavs0_burstcount
	signal mm_interconnect_0_mm_bridge_0_s0_readdata                           : std_logic_vector(31 downto 0); -- mm_bridge_0:s0_readdata -> mm_interconnect_0:mm_bridge_0_s0_readdata
	signal mm_interconnect_0_mm_bridge_0_s0_waitrequest                        : std_logic;                     -- mm_bridge_0:s0_waitrequest -> mm_interconnect_0:mm_bridge_0_s0_waitrequest
	signal mm_interconnect_0_mm_bridge_0_s0_debugaccess                        : std_logic;                     -- mm_interconnect_0:mm_bridge_0_s0_debugaccess -> mm_bridge_0:s0_debugaccess
	signal mm_interconnect_0_mm_bridge_0_s0_address                            : std_logic_vector(14 downto 0); -- mm_interconnect_0:mm_bridge_0_s0_address -> mm_bridge_0:s0_address
	signal mm_interconnect_0_mm_bridge_0_s0_read                               : std_logic;                     -- mm_interconnect_0:mm_bridge_0_s0_read -> mm_bridge_0:s0_read
	signal mm_interconnect_0_mm_bridge_0_s0_byteenable                         : std_logic_vector(3 downto 0);  -- mm_interconnect_0:mm_bridge_0_s0_byteenable -> mm_bridge_0:s0_byteenable
	signal mm_interconnect_0_mm_bridge_0_s0_readdatavalid                      : std_logic;                     -- mm_bridge_0:s0_readdatavalid -> mm_interconnect_0:mm_bridge_0_s0_readdatavalid
	signal mm_interconnect_0_mm_bridge_0_s0_write                              : std_logic;                     -- mm_interconnect_0:mm_bridge_0_s0_write -> mm_bridge_0:s0_write
	signal mm_interconnect_0_mm_bridge_0_s0_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:mm_bridge_0_s0_writedata -> mm_bridge_0:s0_writedata
	signal mm_interconnect_0_mm_bridge_0_s0_burstcount                         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:mm_bridge_0_s0_burstcount -> mm_bridge_0:s0_burstcount
	signal mm_interconnect_0_onchip_ram_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:onchip_ram_s1_chipselect -> onchip_ram:chipselect
	signal mm_interconnect_0_onchip_ram_s1_readdata                            : std_logic_vector(31 downto 0); -- onchip_ram:readdata -> mm_interconnect_0:onchip_ram_s1_readdata
	signal mm_interconnect_0_onchip_ram_s1_address                             : std_logic_vector(8 downto 0);  -- mm_interconnect_0:onchip_ram_s1_address -> onchip_ram:address
	signal mm_interconnect_0_onchip_ram_s1_byteenable                          : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_ram_s1_byteenable -> onchip_ram:byteenable
	signal mm_interconnect_0_onchip_ram_s1_write                               : std_logic;                     -- mm_interconnect_0:onchip_ram_s1_write -> onchip_ram:write
	signal mm_interconnect_0_onchip_ram_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_ram_s1_writedata -> onchip_ram:writedata
	signal mm_interconnect_0_onchip_ram_s1_clken                               : std_logic;                     -- mm_interconnect_0:onchip_ram_s1_clken -> onchip_ram:clken
	signal msgdma_rx_descriptor_read_master_readdata                           : std_logic_vector(31 downto 0); -- mm_interconnect_1:msgdma_rx_descriptor_read_master_readdata -> msgdma_rx:descriptor_read_master_readdata
	signal msgdma_rx_descriptor_read_master_waitrequest                        : std_logic;                     -- mm_interconnect_1:msgdma_rx_descriptor_read_master_waitrequest -> msgdma_rx:descriptor_read_master_waitrequest
	signal msgdma_rx_descriptor_read_master_address                            : std_logic_vector(14 downto 0); -- msgdma_rx:descriptor_read_master_address -> mm_interconnect_1:msgdma_rx_descriptor_read_master_address
	signal msgdma_rx_descriptor_read_master_read                               : std_logic;                     -- msgdma_rx:descriptor_read_master_read -> mm_interconnect_1:msgdma_rx_descriptor_read_master_read
	signal msgdma_rx_descriptor_read_master_readdatavalid                      : std_logic;                     -- mm_interconnect_1:msgdma_rx_descriptor_read_master_readdatavalid -> msgdma_rx:descriptor_read_master_readdatavalid
	signal msgdma_tx_descriptor_read_master_readdata                           : std_logic_vector(31 downto 0); -- mm_interconnect_1:msgdma_tx_descriptor_read_master_readdata -> msgdma_tx:descriptor_read_master_readdata
	signal msgdma_tx_descriptor_read_master_waitrequest                        : std_logic;                     -- mm_interconnect_1:msgdma_tx_descriptor_read_master_waitrequest -> msgdma_tx:descriptor_read_master_waitrequest
	signal msgdma_tx_descriptor_read_master_address                            : std_logic_vector(14 downto 0); -- msgdma_tx:descriptor_read_master_address -> mm_interconnect_1:msgdma_tx_descriptor_read_master_address
	signal msgdma_tx_descriptor_read_master_read                               : std_logic;                     -- msgdma_tx:descriptor_read_master_read -> mm_interconnect_1:msgdma_tx_descriptor_read_master_read
	signal msgdma_tx_descriptor_read_master_readdatavalid                      : std_logic;                     -- mm_interconnect_1:msgdma_tx_descriptor_read_master_readdatavalid -> msgdma_tx:descriptor_read_master_readdatavalid
	signal msgdma_rx_descriptor_write_master_waitrequest                       : std_logic;                     -- mm_interconnect_1:msgdma_rx_descriptor_write_master_waitrequest -> msgdma_rx:descriptor_write_master_waitrequest
	signal msgdma_rx_descriptor_write_master_address                           : std_logic_vector(14 downto 0); -- msgdma_rx:descriptor_write_master_address -> mm_interconnect_1:msgdma_rx_descriptor_write_master_address
	signal msgdma_rx_descriptor_write_master_byteenable                        : std_logic_vector(3 downto 0);  -- msgdma_rx:descriptor_write_master_byteenable -> mm_interconnect_1:msgdma_rx_descriptor_write_master_byteenable
	signal msgdma_rx_descriptor_write_master_response                          : std_logic_vector(1 downto 0);  -- mm_interconnect_1:msgdma_rx_descriptor_write_master_response -> msgdma_rx:descriptor_write_master_response
	signal msgdma_rx_descriptor_write_master_write                             : std_logic;                     -- msgdma_rx:descriptor_write_master_write -> mm_interconnect_1:msgdma_rx_descriptor_write_master_write
	signal msgdma_rx_descriptor_write_master_writedata                         : std_logic_vector(31 downto 0); -- msgdma_rx:descriptor_write_master_writedata -> mm_interconnect_1:msgdma_rx_descriptor_write_master_writedata
	signal msgdma_rx_descriptor_write_master_writeresponsevalid                : std_logic;                     -- mm_interconnect_1:msgdma_rx_descriptor_write_master_writeresponsevalid -> msgdma_rx:descriptor_write_master_writeresponsevalid
	signal msgdma_tx_descriptor_write_master_waitrequest                       : std_logic;                     -- mm_interconnect_1:msgdma_tx_descriptor_write_master_waitrequest -> msgdma_tx:descriptor_write_master_waitrequest
	signal msgdma_tx_descriptor_write_master_address                           : std_logic_vector(14 downto 0); -- msgdma_tx:descriptor_write_master_address -> mm_interconnect_1:msgdma_tx_descriptor_write_master_address
	signal msgdma_tx_descriptor_write_master_byteenable                        : std_logic_vector(3 downto 0);  -- msgdma_tx:descriptor_write_master_byteenable -> mm_interconnect_1:msgdma_tx_descriptor_write_master_byteenable
	signal msgdma_tx_descriptor_write_master_response                          : std_logic_vector(1 downto 0);  -- mm_interconnect_1:msgdma_tx_descriptor_write_master_response -> msgdma_tx:descriptor_write_master_response
	signal msgdma_tx_descriptor_write_master_write                             : std_logic;                     -- msgdma_tx:descriptor_write_master_write -> mm_interconnect_1:msgdma_tx_descriptor_write_master_write
	signal msgdma_tx_descriptor_write_master_writedata                         : std_logic_vector(31 downto 0); -- msgdma_tx:descriptor_write_master_writedata -> mm_interconnect_1:msgdma_tx_descriptor_write_master_writedata
	signal msgdma_tx_descriptor_write_master_writeresponsevalid                : std_logic;                     -- mm_interconnect_1:msgdma_tx_descriptor_write_master_writeresponsevalid -> msgdma_tx:descriptor_write_master_writeresponsevalid
	signal mm_bridge_0_m0_waitrequest                                          : std_logic;                     -- mm_interconnect_1:mm_bridge_0_m0_waitrequest -> mm_bridge_0:m0_waitrequest
	signal mm_bridge_0_m0_readdata                                             : std_logic_vector(31 downto 0); -- mm_interconnect_1:mm_bridge_0_m0_readdata -> mm_bridge_0:m0_readdata
	signal mm_bridge_0_m0_debugaccess                                          : std_logic;                     -- mm_bridge_0:m0_debugaccess -> mm_interconnect_1:mm_bridge_0_m0_debugaccess
	signal mm_bridge_0_m0_address                                              : std_logic_vector(14 downto 0); -- mm_bridge_0:m0_address -> mm_interconnect_1:mm_bridge_0_m0_address
	signal mm_bridge_0_m0_read                                                 : std_logic;                     -- mm_bridge_0:m0_read -> mm_interconnect_1:mm_bridge_0_m0_read
	signal mm_bridge_0_m0_byteenable                                           : std_logic_vector(3 downto 0);  -- mm_bridge_0:m0_byteenable -> mm_interconnect_1:mm_bridge_0_m0_byteenable
	signal mm_bridge_0_m0_readdatavalid                                        : std_logic;                     -- mm_interconnect_1:mm_bridge_0_m0_readdatavalid -> mm_bridge_0:m0_readdatavalid
	signal mm_bridge_0_m0_writedata                                            : std_logic_vector(31 downto 0); -- mm_bridge_0:m0_writedata -> mm_interconnect_1:mm_bridge_0_m0_writedata
	signal mm_bridge_0_m0_write                                                : std_logic;                     -- mm_bridge_0:m0_write -> mm_interconnect_1:mm_bridge_0_m0_write
	signal mm_bridge_0_m0_burstcount                                           : std_logic_vector(0 downto 0);  -- mm_bridge_0:m0_burstcount -> mm_interconnect_1:mm_bridge_0_m0_burstcount
	signal mm_interconnect_1_descriptor_memory_s1_chipselect                   : std_logic;                     -- mm_interconnect_1:descriptor_memory_s1_chipselect -> descriptor_memory:chipselect
	signal mm_interconnect_1_descriptor_memory_s1_readdata                     : std_logic_vector(31 downto 0); -- descriptor_memory:readdata -> mm_interconnect_1:descriptor_memory_s1_readdata
	signal mm_interconnect_1_descriptor_memory_s1_address                      : std_logic_vector(10 downto 0); -- mm_interconnect_1:descriptor_memory_s1_address -> descriptor_memory:address
	signal mm_interconnect_1_descriptor_memory_s1_byteenable                   : std_logic_vector(3 downto 0);  -- mm_interconnect_1:descriptor_memory_s1_byteenable -> descriptor_memory:byteenable
	signal mm_interconnect_1_descriptor_memory_s1_write                        : std_logic;                     -- mm_interconnect_1:descriptor_memory_s1_write -> descriptor_memory:write
	signal mm_interconnect_1_descriptor_memory_s1_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_1:descriptor_memory_s1_writedata -> descriptor_memory:writedata
	signal mm_interconnect_1_descriptor_memory_s1_clken                        : std_logic;                     -- mm_interconnect_1:descriptor_memory_s1_clken -> descriptor_memory:clken
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect            : std_logic;                     -- mm_interconnect_1:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata              : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest           : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_address               : std_logic_vector(0 downto 0);  -- mm_interconnect_1:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_read                  : std_logic;                     -- mm_interconnect_1:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_1_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_write                 : std_logic;                     -- mm_interconnect_1:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_1_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_1:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_1_opencores_i2c_0_avalon_slave_0_chipselect         : std_logic;                     -- mm_interconnect_1:opencores_i2c_0_avalon_slave_0_chipselect -> opencores_i2c_0:wb_stb_i
	signal mm_interconnect_1_opencores_i2c_0_avalon_slave_0_readdata           : std_logic_vector(7 downto 0);  -- opencores_i2c_0:wb_dat_o -> mm_interconnect_1:opencores_i2c_0_avalon_slave_0_readdata
	signal opencores_i2c_0_avalon_slave_0_waitrequest                          : std_logic;                     -- opencores_i2c_0:wb_ack_o -> opencores_i2c_0_avalon_slave_0_waitrequest:in
	signal mm_interconnect_1_opencores_i2c_0_avalon_slave_0_address            : std_logic_vector(2 downto 0);  -- mm_interconnect_1:opencores_i2c_0_avalon_slave_0_address -> opencores_i2c_0:wb_adr_i
	signal mm_interconnect_1_opencores_i2c_0_avalon_slave_0_write              : std_logic;                     -- mm_interconnect_1:opencores_i2c_0_avalon_slave_0_write -> opencores_i2c_0:wb_we_i
	signal mm_interconnect_1_opencores_i2c_0_avalon_slave_0_writedata          : std_logic_vector(7 downto 0);  -- mm_interconnect_1:opencores_i2c_0_avalon_slave_0_writedata -> opencores_i2c_0:wb_dat_i
	signal mm_interconnect_1_userhw_0_avalon_slave_0_readdata                  : std_logic_vector(31 downto 0); -- userhw_0:readdata -> mm_interconnect_1:userhw_0_avalon_slave_0_readdata
	signal mm_interconnect_1_userhw_0_avalon_slave_0_address                   : std_logic_vector(2 downto 0);  -- mm_interconnect_1:userhw_0_avalon_slave_0_address -> userhw_0:address
	signal mm_interconnect_1_userhw_0_avalon_slave_0_read                      : std_logic;                     -- mm_interconnect_1:userhw_0_avalon_slave_0_read -> userhw_0:read
	signal mm_interconnect_1_userhw_0_avalon_slave_0_write                     : std_logic;                     -- mm_interconnect_1:userhw_0_avalon_slave_0_write -> userhw_0:write
	signal mm_interconnect_1_userhw_0_avalon_slave_0_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_1:userhw_0_avalon_slave_0_writedata -> userhw_0:writedata
	signal mm_interconnect_1_eth_tse_control_port_readdata                     : std_logic_vector(31 downto 0); -- eth_tse:reg_data_out -> mm_interconnect_1:eth_tse_control_port_readdata
	signal mm_interconnect_1_eth_tse_control_port_waitrequest                  : std_logic;                     -- eth_tse:reg_busy -> mm_interconnect_1:eth_tse_control_port_waitrequest
	signal mm_interconnect_1_eth_tse_control_port_address                      : std_logic_vector(7 downto 0);  -- mm_interconnect_1:eth_tse_control_port_address -> eth_tse:reg_addr
	signal mm_interconnect_1_eth_tse_control_port_read                         : std_logic;                     -- mm_interconnect_1:eth_tse_control_port_read -> eth_tse:reg_rd
	signal mm_interconnect_1_eth_tse_control_port_write                        : std_logic;                     -- mm_interconnect_1:eth_tse_control_port_write -> eth_tse:reg_wr
	signal mm_interconnect_1_eth_tse_control_port_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_1:eth_tse_control_port_writedata -> eth_tse:reg_data_in
	signal mm_interconnect_1_sysid_control_slave_readdata                      : std_logic_vector(31 downto 0); -- sysid:readdata -> mm_interconnect_1:sysid_control_slave_readdata
	signal mm_interconnect_1_sysid_control_slave_address                       : std_logic_vector(0 downto 0);  -- mm_interconnect_1:sysid_control_slave_address -> sysid:address
	signal mm_interconnect_1_msgdma_rx_csr_readdata                            : std_logic_vector(31 downto 0); -- msgdma_rx:csr_readdata -> mm_interconnect_1:msgdma_rx_csr_readdata
	signal mm_interconnect_1_msgdma_rx_csr_address                             : std_logic_vector(2 downto 0);  -- mm_interconnect_1:msgdma_rx_csr_address -> msgdma_rx:csr_address
	signal mm_interconnect_1_msgdma_rx_csr_read                                : std_logic;                     -- mm_interconnect_1:msgdma_rx_csr_read -> msgdma_rx:csr_read
	signal mm_interconnect_1_msgdma_rx_csr_byteenable                          : std_logic_vector(3 downto 0);  -- mm_interconnect_1:msgdma_rx_csr_byteenable -> msgdma_rx:csr_byteenable
	signal mm_interconnect_1_msgdma_rx_csr_write                               : std_logic;                     -- mm_interconnect_1:msgdma_rx_csr_write -> msgdma_rx:csr_write
	signal mm_interconnect_1_msgdma_rx_csr_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_1:msgdma_rx_csr_writedata -> msgdma_rx:csr_writedata
	signal mm_interconnect_1_msgdma_tx_csr_readdata                            : std_logic_vector(31 downto 0); -- msgdma_tx:csr_readdata -> mm_interconnect_1:msgdma_tx_csr_readdata
	signal mm_interconnect_1_msgdma_tx_csr_address                             : std_logic_vector(2 downto 0);  -- mm_interconnect_1:msgdma_tx_csr_address -> msgdma_tx:csr_address
	signal mm_interconnect_1_msgdma_tx_csr_read                                : std_logic;                     -- mm_interconnect_1:msgdma_tx_csr_read -> msgdma_tx:csr_read
	signal mm_interconnect_1_msgdma_tx_csr_byteenable                          : std_logic_vector(3 downto 0);  -- mm_interconnect_1:msgdma_tx_csr_byteenable -> msgdma_tx:csr_byteenable
	signal mm_interconnect_1_msgdma_tx_csr_write                               : std_logic;                     -- mm_interconnect_1:msgdma_tx_csr_write -> msgdma_tx:csr_write
	signal mm_interconnect_1_msgdma_tx_csr_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_1:msgdma_tx_csr_writedata -> msgdma_tx:csr_writedata
	signal mm_interconnect_1_msgdma_tx_prefetcher_csr_readdata                 : std_logic_vector(31 downto 0); -- msgdma_tx:prefetcher_csr_readdata -> mm_interconnect_1:msgdma_tx_prefetcher_csr_readdata
	signal mm_interconnect_1_msgdma_tx_prefetcher_csr_address                  : std_logic_vector(2 downto 0);  -- mm_interconnect_1:msgdma_tx_prefetcher_csr_address -> msgdma_tx:prefetcher_csr_address
	signal mm_interconnect_1_msgdma_tx_prefetcher_csr_read                     : std_logic;                     -- mm_interconnect_1:msgdma_tx_prefetcher_csr_read -> msgdma_tx:prefetcher_csr_read
	signal mm_interconnect_1_msgdma_tx_prefetcher_csr_write                    : std_logic;                     -- mm_interconnect_1:msgdma_tx_prefetcher_csr_write -> msgdma_tx:prefetcher_csr_write
	signal mm_interconnect_1_msgdma_tx_prefetcher_csr_writedata                : std_logic_vector(31 downto 0); -- mm_interconnect_1:msgdma_tx_prefetcher_csr_writedata -> msgdma_tx:prefetcher_csr_writedata
	signal mm_interconnect_1_msgdma_rx_prefetcher_csr_readdata                 : std_logic_vector(31 downto 0); -- msgdma_rx:prefetcher_csr_readdata -> mm_interconnect_1:msgdma_rx_prefetcher_csr_readdata
	signal mm_interconnect_1_msgdma_rx_prefetcher_csr_address                  : std_logic_vector(2 downto 0);  -- mm_interconnect_1:msgdma_rx_prefetcher_csr_address -> msgdma_rx:prefetcher_csr_address
	signal mm_interconnect_1_msgdma_rx_prefetcher_csr_read                     : std_logic;                     -- mm_interconnect_1:msgdma_rx_prefetcher_csr_read -> msgdma_rx:prefetcher_csr_read
	signal mm_interconnect_1_msgdma_rx_prefetcher_csr_write                    : std_logic;                     -- mm_interconnect_1:msgdma_rx_prefetcher_csr_write -> msgdma_rx:prefetcher_csr_write
	signal mm_interconnect_1_msgdma_rx_prefetcher_csr_writedata                : std_logic_vector(31 downto 0); -- mm_interconnect_1:msgdma_rx_prefetcher_csr_writedata -> msgdma_rx:prefetcher_csr_writedata
	signal mm_interconnect_1_sys_clk_timer_s1_chipselect                       : std_logic;                     -- mm_interconnect_1:sys_clk_timer_s1_chipselect -> sys_clk_timer:chipselect
	signal mm_interconnect_1_sys_clk_timer_s1_readdata                         : std_logic_vector(15 downto 0); -- sys_clk_timer:readdata -> mm_interconnect_1:sys_clk_timer_s1_readdata
	signal mm_interconnect_1_sys_clk_timer_s1_address                          : std_logic_vector(2 downto 0);  -- mm_interconnect_1:sys_clk_timer_s1_address -> sys_clk_timer:address
	signal mm_interconnect_1_sys_clk_timer_s1_write                            : std_logic;                     -- mm_interconnect_1:sys_clk_timer_s1_write -> mm_interconnect_1_sys_clk_timer_s1_write:in
	signal mm_interconnect_1_sys_clk_timer_s1_writedata                        : std_logic_vector(15 downto 0); -- mm_interconnect_1:sys_clk_timer_s1_writedata -> sys_clk_timer:writedata
	signal mm_interconnect_1_led_pio_s1_chipselect                             : std_logic;                     -- mm_interconnect_1:led_pio_s1_chipselect -> led_pio:chipselect
	signal mm_interconnect_1_led_pio_s1_readdata                               : std_logic_vector(31 downto 0); -- led_pio:readdata -> mm_interconnect_1:led_pio_s1_readdata
	signal mm_interconnect_1_led_pio_s1_address                                : std_logic_vector(1 downto 0);  -- mm_interconnect_1:led_pio_s1_address -> led_pio:address
	signal mm_interconnect_1_led_pio_s1_write                                  : std_logic;                     -- mm_interconnect_1:led_pio_s1_write -> mm_interconnect_1_led_pio_s1_write:in
	signal mm_interconnect_1_led_pio_s1_writedata                              : std_logic_vector(31 downto 0); -- mm_interconnect_1:led_pio_s1_writedata -> led_pio:writedata
	signal mm_interconnect_1_user_dipsw_s1_readdata                            : std_logic_vector(31 downto 0); -- user_dipsw:readdata -> mm_interconnect_1:user_dipsw_s1_readdata
	signal mm_interconnect_1_user_dipsw_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_1:user_dipsw_s1_address -> user_dipsw:address
	signal mm_interconnect_1_user_pb_s1_readdata                               : std_logic_vector(31 downto 0); -- user_pb:readdata -> mm_interconnect_1:user_pb_s1_readdata
	signal mm_interconnect_1_user_pb_s1_address                                : std_logic_vector(1 downto 0);  -- mm_interconnect_1:user_pb_s1_address -> user_pb:address
	signal irq_mapper_receiver0_irq                                            : std_logic;                     -- msgdma_rx:csr_irq_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                            : std_logic;                     -- msgdma_tx:csr_irq_irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                            : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                            : std_logic;                     -- sys_clk_timer:irq -> irq_mapper:receiver3_irq
	signal cpu_irq_irq                                                         : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> cpu:irq
	signal eth_tse_receive_valid                                               : std_logic;                     -- eth_tse:ff_rx_dval -> avalon_st_adapter:in_0_valid
	signal eth_tse_receive_data                                                : std_logic_vector(31 downto 0); -- eth_tse:ff_rx_data -> avalon_st_adapter:in_0_data
	signal eth_tse_receive_ready                                               : std_logic;                     -- avalon_st_adapter:in_0_ready -> eth_tse:ff_rx_rdy
	signal eth_tse_receive_startofpacket                                       : std_logic;                     -- eth_tse:ff_rx_sop -> avalon_st_adapter:in_0_startofpacket
	signal eth_tse_receive_endofpacket                                         : std_logic;                     -- eth_tse:ff_rx_eop -> avalon_st_adapter:in_0_endofpacket
	signal eth_tse_receive_error                                               : std_logic_vector(5 downto 0);  -- eth_tse:rx_err -> avalon_st_adapter:in_0_error
	signal eth_tse_receive_empty                                               : std_logic_vector(1 downto 0);  -- eth_tse:ff_rx_mod -> avalon_st_adapter:in_0_empty
	signal avalon_st_adapter_out_0_valid                                       : std_logic;                     -- avalon_st_adapter:out_0_valid -> msgdma_rx:st_sink_valid
	signal avalon_st_adapter_out_0_data                                        : std_logic_vector(31 downto 0); -- avalon_st_adapter:out_0_data -> msgdma_rx:st_sink_data
	signal avalon_st_adapter_out_0_ready                                       : std_logic;                     -- msgdma_rx:st_sink_ready -> avalon_st_adapter:out_0_ready
	signal avalon_st_adapter_out_0_startofpacket                               : std_logic;                     -- avalon_st_adapter:out_0_startofpacket -> msgdma_rx:st_sink_startofpacket
	signal avalon_st_adapter_out_0_endofpacket                                 : std_logic;                     -- avalon_st_adapter:out_0_endofpacket -> msgdma_rx:st_sink_endofpacket
	signal avalon_st_adapter_out_0_error                                       : std_logic_vector(5 downto 0);  -- avalon_st_adapter:out_0_error -> msgdma_rx:st_sink_error
	signal avalon_st_adapter_out_0_empty                                       : std_logic_vector(1 downto 0);  -- avalon_st_adapter:out_0_empty -> msgdma_rx:st_sink_empty
	signal rst_controller_reset_out_reset                                      : std_logic;                     -- rst_controller:reset_out -> [avalon_st_adapter:in_rst_0_reset, descriptor_memory:reset, eth_tse:reset, irq_mapper:reset, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, mm_interconnect_1:descriptor_memory_reset1_reset_bridge_in_reset_reset, onchip_ram:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                                  : std_logic;                     -- rst_controller:reset_req -> [cpu:reset_req, descriptor_memory:reset_req, onchip_ram:reset_req, rst_translator:reset_req_in]
	signal cpu_debug_reset_request_reset                                       : std_logic;                     -- cpu:debug_reset_request -> rst_controller:reset_in0
	signal rst_controller_001_reset_out_reset                                  : std_logic;                     -- rst_controller_001:reset_out -> enet_pll:reset
	signal rst_controller_002_reset_out_reset                                  : std_logic;                     -- rst_controller_002:reset_out -> [mm_interconnect_0:ext_epcq_flash_reset_reset_bridge_in_reset_reset, remote_update:reset_reset, rst_controller_002_reset_out_reset:in]
	signal rst_controller_003_reset_out_reset                                  : std_logic;                     -- rst_controller_003:reset_out -> rst_controller_003_reset_out_reset:in
	signal hbus_reset_reset_n_ports_inv                                        : std_logic;                     -- hbus_reset_reset_n:inv -> [rst_controller_002:reset_in0, rst_controller_003:reset_in0]
	signal reset_enet_reset_n_ports_inv                                        : std_logic;                     -- reset_enet_reset_n:inv -> rst_controller_001:reset_in0
	signal sll_hyperbus_controller_top_0_o_av_out_rstn_reset_ports_inv         : std_logic;                     -- sll_hyperbus_controller_top_0_o_av_out_rstn_reset:inv -> [mm_bridge_0:reset, mm_interconnect_0:sll_hyperbus_controller_top_0_i_iavs0_rstn_reset_bridge_in_reset_reset, mm_interconnect_1:msgdma_rx_reset_n_reset_bridge_in_reset_reset, opencores_i2c_0:wb_rst_i, rst_controller:reset_in1, userhw_0:rst]
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_read_ports_inv        : std_logic;                     -- mm_interconnect_1_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_write_ports_inv       : std_logic;                     -- mm_interconnect_1_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_1_opencores_i2c_0_avalon_slave_0_inv                : std_logic;                     -- opencores_i2c_0_avalon_slave_0_waitrequest:inv -> mm_interconnect_1:opencores_i2c_0_avalon_slave_0_waitrequest
	signal mm_interconnect_1_sys_clk_timer_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_1_sys_clk_timer_s1_write:inv -> sys_clk_timer:write_n
	signal mm_interconnect_1_led_pio_s1_write_ports_inv                        : std_logic;                     -- mm_interconnect_1_led_pio_s1_write:inv -> led_pio:write_n
	signal rst_controller_reset_out_reset_ports_inv                            : std_logic;                     -- rst_controller_reset_out_reset:inv -> [cpu:reset_n, jtag_uart:rst_n, led_pio:reset_n, sys_clk_timer:reset_n, sysid:reset_n]
	signal rst_controller_002_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_002_reset_out_reset:inv -> ext_epcq_flash:reset_n
	signal rst_controller_003_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_003_reset_out_reset:inv -> sll_hyperbus_controller_top_0:i_ext_rstn

begin

	cpu : component q_sys_cpu
		port map (
			clk                                 => sll_hyperbus_controller_top_0_o_av_out_clk_clk,    --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,          --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                --                          .reset_req
			d_address                           => cpu_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_data_master_read,                              --                          .read
			d_readdata                          => cpu_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_data_master_write,                             --                          .write
			d_writedata                         => cpu_data_master_writedata,                         --                          .writedata
			d_burstcount                        => cpu_data_master_burstcount,                        --                          .burstcount
			d_readdatavalid                     => cpu_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => cpu_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_instruction_master_waitrequest,                --                          .waitrequest
			i_burstcount                        => cpu_instruction_master_burstcount,                 --                          .burstcount
			i_readdatavalid                     => cpu_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => cpu_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => cpu_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                               -- custom_instruction_master.readra
		);

	descriptor_memory : component q_sys_descriptor_memory
		port map (
			clk        => sll_hyperbus_controller_top_0_o_av_out_clk_clk,    --   clk1.clk
			address    => mm_interconnect_1_descriptor_memory_s1_address,    --     s1.address
			clken      => mm_interconnect_1_descriptor_memory_s1_clken,      --       .clken
			chipselect => mm_interconnect_1_descriptor_memory_s1_chipselect, --       .chipselect
			write      => mm_interconnect_1_descriptor_memory_s1_write,      --       .write
			readdata   => mm_interconnect_1_descriptor_memory_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_1_descriptor_memory_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_1_descriptor_memory_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                    -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,                --       .reset_req
			freeze     => '0'                                                -- (terminated)
		);

	enet_pll : component q_sys_enet_pll
		port map (
			clk                => enet_clk_125m_in_clk,               --       inclk_interface.clk
			reset              => rst_controller_001_reset_out_reset, -- inclk_interface_reset.reset
			read               => open,                               --             pll_slave.read
			write              => open,                               --                      .write
			address            => open,                               --                      .address
			readdata           => open,                               --                      .readdata
			writedata          => open,                               --                      .writedata
			c0                 => enet_pll_c0_125m_clk,               --                    c0.clk
			c1                 => enet_pll_c1_25m_clk,                --                    c1.clk
			c2                 => enet_pll_c2_2m5_clk,                --                    c2.clk
			c3                 => enet_pll_c3_125m_shift_clk,         --                    c3.clk
			c4                 => enet_pll_c4_25m_shift_clk,          --                    c4.clk
			areset             => enet_pll_areset_conduit_export,     --        areset_conduit.export
			locked             => enet_pll_locked_conduit_export,     --        locked_conduit.export
			scandone           => open,                               --           (terminated)
			scandataout        => open,                               --           (terminated)
			phasedone          => open,                               --           (terminated)
			phasecounterselect => "0000",                             --           (terminated)
			phaseupdown        => '0',                                --           (terminated)
			phasestep          => '0',                                --           (terminated)
			scanclk            => '0',                                --           (terminated)
			scanclkena         => '0',                                --           (terminated)
			scandata           => '0',                                --           (terminated)
			configupdate       => '0'                                 --           (terminated)
		);

	eth_tse : component q_sys_eth_tse
		port map (
			clk           => sll_hyperbus_controller_top_0_o_av_out_clk_clk,     -- control_port_clock_connection.clk
			reset         => rst_controller_reset_out_reset,                     --              reset_connection.reset
			reg_addr      => mm_interconnect_1_eth_tse_control_port_address,     --                  control_port.address
			reg_data_out  => mm_interconnect_1_eth_tse_control_port_readdata,    --                              .readdata
			reg_rd        => mm_interconnect_1_eth_tse_control_port_read,        --                              .read
			reg_data_in   => mm_interconnect_1_eth_tse_control_port_writedata,   --                              .writedata
			reg_wr        => mm_interconnect_1_eth_tse_control_port_write,       --                              .write
			reg_busy      => mm_interconnect_1_eth_tse_control_port_waitrequest, --                              .waitrequest
			tx_clk        => eth_tse_pcs_mac_tx_clock_connection_clk,            --   pcs_mac_tx_clock_connection.clk
			rx_clk        => eth_tse_pcs_mac_rx_clock_connection_clk,            --   pcs_mac_rx_clock_connection.clk
			set_10        => eth_tse_mac_status_connection_set_10,               --         mac_status_connection.set_10
			set_1000      => eth_tse_mac_status_connection_set_1000,             --                              .set_1000
			eth_mode      => eth_tse_mac_status_connection_eth_mode,             --                              .eth_mode
			ena_10        => eth_tse_mac_status_connection_ena_10,               --                              .ena_10
			rgmii_in      => eth_tse_mac_rgmii_connection_rgmii_in,              --          mac_rgmii_connection.rgmii_in
			rgmii_out     => eth_tse_mac_rgmii_connection_rgmii_out,             --                              .rgmii_out
			rx_control    => eth_tse_mac_rgmii_connection_rx_control,            --                              .rx_control
			tx_control    => eth_tse_mac_rgmii_connection_tx_control,            --                              .tx_control
			ff_rx_clk     => sll_hyperbus_controller_top_0_o_av_out_clk_clk,     --      receive_clock_connection.clk
			ff_tx_clk     => sll_hyperbus_controller_top_0_o_av_out_clk_clk,     --     transmit_clock_connection.clk
			ff_rx_data    => eth_tse_receive_data,                               --                       receive.data
			ff_rx_eop     => eth_tse_receive_endofpacket,                        --                              .endofpacket
			rx_err        => eth_tse_receive_error,                              --                              .error
			ff_rx_mod     => eth_tse_receive_empty,                              --                              .empty
			ff_rx_rdy     => eth_tse_receive_ready,                              --                              .ready
			ff_rx_sop     => eth_tse_receive_startofpacket,                      --                              .startofpacket
			ff_rx_dval    => eth_tse_receive_valid,                              --                              .valid
			ff_tx_data    => msgdma_tx_st_source_data,                           --                      transmit.data
			ff_tx_eop     => msgdma_tx_st_source_endofpacket,                    --                              .endofpacket
			ff_tx_err     => msgdma_tx_st_source_error,                          --                              .error
			ff_tx_mod     => msgdma_tx_st_source_empty,                          --                              .empty
			ff_tx_rdy     => msgdma_tx_st_source_ready,                          --                              .ready
			ff_tx_sop     => msgdma_tx_st_source_startofpacket,                  --                              .startofpacket
			ff_tx_wren    => msgdma_tx_st_source_valid,                          --                              .valid
			mdc           => eth_tse_mac_mdio_connection_mdc,                    --           mac_mdio_connection.mdc
			mdio_in       => eth_tse_mac_mdio_connection_mdio_in,                --                              .mdio_in
			mdio_out      => eth_tse_mac_mdio_connection_mdio_out,               --                              .mdio_out
			mdio_oen      => eth_tse_mac_mdio_connection_mdio_oen,               --                              .mdio_oen
			magic_wakeup  => open,                                               --           mac_misc_connection.magic_wakeup
			magic_sleep_n => open,                                               --                              .magic_sleep_n
			ff_tx_crc_fwd => open,                                               --                              .ff_tx_crc_fwd
			ff_tx_septy   => open,                                               --                              .ff_tx_septy
			tx_ff_uflow   => open,                                               --                              .tx_ff_uflow
			ff_tx_a_full  => open,                                               --                              .ff_tx_a_full
			ff_tx_a_empty => open,                                               --                              .ff_tx_a_empty
			rx_err_stat   => open,                                               --                              .rx_err_stat
			rx_frm_type   => open,                                               --                              .rx_frm_type
			ff_rx_dsav    => open,                                               --                              .ff_rx_dsav
			ff_rx_a_full  => open,                                               --                              .ff_rx_a_full
			ff_rx_a_empty => open                                                --                              .ff_rx_a_empty
		);

	ext_epcq_flash : component q_sys_ext_epcq_flash
		generic map (
			DEVICE_FAMILY     => "Cyclone 10 LP",
			ASI_WIDTH         => 1,
			CS_WIDTH          => 1,
			ADDR_WIDTH        => 21,
			ASMI_ADDR_WIDTH   => 24,
			ENABLE_4BYTE_ADDR => 0,
			CHIP_SELS         => 1
		)
		port map (
			avl_csr_read         => mm_interconnect_0_ext_epcq_flash_avl_csr_read,          --          avl_csr.read
			avl_csr_waitrequest  => mm_interconnect_0_ext_epcq_flash_avl_csr_waitrequest,   --                 .waitrequest
			avl_csr_write        => mm_interconnect_0_ext_epcq_flash_avl_csr_write,         --                 .write
			avl_csr_addr         => mm_interconnect_0_ext_epcq_flash_avl_csr_address,       --                 .address
			avl_csr_wrdata       => mm_interconnect_0_ext_epcq_flash_avl_csr_writedata,     --                 .writedata
			avl_csr_rddata       => mm_interconnect_0_ext_epcq_flash_avl_csr_readdata,      --                 .readdata
			avl_csr_rddata_valid => mm_interconnect_0_ext_epcq_flash_avl_csr_readdatavalid, --                 .readdatavalid
			avl_mem_write        => mm_interconnect_0_ext_epcq_flash_avl_mem_write,         --          avl_mem.write
			avl_mem_burstcount   => mm_interconnect_0_ext_epcq_flash_avl_mem_burstcount,    --                 .burstcount
			avl_mem_waitrequest  => mm_interconnect_0_ext_epcq_flash_avl_mem_waitrequest,   --                 .waitrequest
			avl_mem_read         => mm_interconnect_0_ext_epcq_flash_avl_mem_read,          --                 .read
			avl_mem_addr         => mm_interconnect_0_ext_epcq_flash_avl_mem_address,       --                 .address
			avl_mem_wrdata       => mm_interconnect_0_ext_epcq_flash_avl_mem_writedata,     --                 .writedata
			avl_mem_rddata       => mm_interconnect_0_ext_epcq_flash_avl_mem_readdata,      --                 .readdata
			avl_mem_rddata_valid => mm_interconnect_0_ext_epcq_flash_avl_mem_readdatavalid, --                 .readdatavalid
			avl_mem_byteenable   => mm_interconnect_0_ext_epcq_flash_avl_mem_byteenable,    --                 .byteenable
			irq                  => open,                                                   -- interrupt_sender.irq
			clk                  => clock_bridge_0_in_clk_clk,                              --       clock_sink.clk
			reset_n              => rst_controller_002_reset_out_reset_ports_inv            --            reset.reset_n
		);

	jtag_uart : component q_sys_jtag_uart
		port map (
			clk            => sll_hyperbus_controller_top_0_o_av_out_clk_clk,                --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_1_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_1_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_1_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver2_irq                                       --               irq.irq
		);

	led_pio : component q_sys_led_pio
		port map (
			clk        => sll_hyperbus_controller_top_0_o_av_out_clk_clk, --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,       --               reset.reset_n
			address    => mm_interconnect_1_led_pio_s1_address,           --                  s1.address
			write_n    => mm_interconnect_1_led_pio_s1_write_ports_inv,   --                    .write_n
			writedata  => mm_interconnect_1_led_pio_s1_writedata,         --                    .writedata
			chipselect => mm_interconnect_1_led_pio_s1_chipselect,        --                    .chipselect
			readdata   => mm_interconnect_1_led_pio_s1_readdata,          --                    .readdata
			out_port   => led_pio_external_connection_export              -- external_connection.export
		);

	mm_bridge_0 : component altera_avalon_mm_bridge
		generic map (
			DATA_WIDTH        => 32,
			SYMBOL_WIDTH      => 8,
			HDL_ADDR_WIDTH    => 15,
			BURSTCOUNT_WIDTH  => 1,
			PIPELINE_COMMAND  => 1,
			PIPELINE_RESPONSE => 1
		)
		port map (
			clk              => sll_hyperbus_controller_top_0_o_av_out_clk_clk,              --   clk.clk
			reset            => sll_hyperbus_controller_top_0_o_av_out_rstn_reset_ports_inv, -- reset.reset
			s0_waitrequest   => mm_interconnect_0_mm_bridge_0_s0_waitrequest,                --    s0.waitrequest
			s0_readdata      => mm_interconnect_0_mm_bridge_0_s0_readdata,                   --      .readdata
			s0_readdatavalid => mm_interconnect_0_mm_bridge_0_s0_readdatavalid,              --      .readdatavalid
			s0_burstcount    => mm_interconnect_0_mm_bridge_0_s0_burstcount,                 --      .burstcount
			s0_writedata     => mm_interconnect_0_mm_bridge_0_s0_writedata,                  --      .writedata
			s0_address       => mm_interconnect_0_mm_bridge_0_s0_address,                    --      .address
			s0_write         => mm_interconnect_0_mm_bridge_0_s0_write,                      --      .write
			s0_read          => mm_interconnect_0_mm_bridge_0_s0_read,                       --      .read
			s0_byteenable    => mm_interconnect_0_mm_bridge_0_s0_byteenable,                 --      .byteenable
			s0_debugaccess   => mm_interconnect_0_mm_bridge_0_s0_debugaccess,                --      .debugaccess
			m0_waitrequest   => mm_bridge_0_m0_waitrequest,                                  --    m0.waitrequest
			m0_readdata      => mm_bridge_0_m0_readdata,                                     --      .readdata
			m0_readdatavalid => mm_bridge_0_m0_readdatavalid,                                --      .readdatavalid
			m0_burstcount    => mm_bridge_0_m0_burstcount,                                   --      .burstcount
			m0_writedata     => mm_bridge_0_m0_writedata,                                    --      .writedata
			m0_address       => mm_bridge_0_m0_address,                                      --      .address
			m0_write         => mm_bridge_0_m0_write,                                        --      .write
			m0_read          => mm_bridge_0_m0_read,                                         --      .read
			m0_byteenable    => mm_bridge_0_m0_byteenable,                                   --      .byteenable
			m0_debugaccess   => mm_bridge_0_m0_debugaccess,                                  --      .debugaccess
			s0_response      => open,                                                        -- (terminated)
			m0_response      => "00"                                                         -- (terminated)
		);

	msgdma_rx : component q_sys_msgdma_rx
		port map (
			mm_write_address                           => msgdma_rx_mm_write_address,                           --                mm_write.address
			mm_write_write                             => msgdma_rx_mm_write_write,                             --                        .write
			mm_write_byteenable                        => msgdma_rx_mm_write_byteenable,                        --                        .byteenable
			mm_write_writedata                         => msgdma_rx_mm_write_writedata,                         --                        .writedata
			mm_write_waitrequest                       => msgdma_rx_mm_write_waitrequest,                       --                        .waitrequest
			descriptor_read_master_address             => msgdma_rx_descriptor_read_master_address,             --  descriptor_read_master.address
			descriptor_read_master_read                => msgdma_rx_descriptor_read_master_read,                --                        .read
			descriptor_read_master_readdata            => msgdma_rx_descriptor_read_master_readdata,            --                        .readdata
			descriptor_read_master_waitrequest         => msgdma_rx_descriptor_read_master_waitrequest,         --                        .waitrequest
			descriptor_read_master_readdatavalid       => msgdma_rx_descriptor_read_master_readdatavalid,       --                        .readdatavalid
			descriptor_write_master_address            => msgdma_rx_descriptor_write_master_address,            -- descriptor_write_master.address
			descriptor_write_master_write              => msgdma_rx_descriptor_write_master_write,              --                        .write
			descriptor_write_master_byteenable         => msgdma_rx_descriptor_write_master_byteenable,         --                        .byteenable
			descriptor_write_master_writedata          => msgdma_rx_descriptor_write_master_writedata,          --                        .writedata
			descriptor_write_master_waitrequest        => msgdma_rx_descriptor_write_master_waitrequest,        --                        .waitrequest
			descriptor_write_master_response           => msgdma_rx_descriptor_write_master_response,           --                        .response
			descriptor_write_master_writeresponsevalid => msgdma_rx_descriptor_write_master_writeresponsevalid, --                        .writeresponsevalid
			clock_clk                                  => sll_hyperbus_controller_top_0_o_av_out_clk_clk,       --                   clock.clk
			reset_n_reset_n                            => sll_hyperbus_controller_top_0_o_av_out_rstn_reset,    --                 reset_n.reset_n
			csr_writedata                              => mm_interconnect_1_msgdma_rx_csr_writedata,            --                     csr.writedata
			csr_write                                  => mm_interconnect_1_msgdma_rx_csr_write,                --                        .write
			csr_byteenable                             => mm_interconnect_1_msgdma_rx_csr_byteenable,           --                        .byteenable
			csr_readdata                               => mm_interconnect_1_msgdma_rx_csr_readdata,             --                        .readdata
			csr_read                                   => mm_interconnect_1_msgdma_rx_csr_read,                 --                        .read
			csr_address                                => mm_interconnect_1_msgdma_rx_csr_address,              --                        .address
			prefetcher_csr_address                     => mm_interconnect_1_msgdma_rx_prefetcher_csr_address,   --          prefetcher_csr.address
			prefetcher_csr_read                        => mm_interconnect_1_msgdma_rx_prefetcher_csr_read,      --                        .read
			prefetcher_csr_write                       => mm_interconnect_1_msgdma_rx_prefetcher_csr_write,     --                        .write
			prefetcher_csr_writedata                   => mm_interconnect_1_msgdma_rx_prefetcher_csr_writedata, --                        .writedata
			prefetcher_csr_readdata                    => mm_interconnect_1_msgdma_rx_prefetcher_csr_readdata,  --                        .readdata
			csr_irq_irq                                => irq_mapper_receiver0_irq,                             --                 csr_irq.irq
			st_sink_data                               => avalon_st_adapter_out_0_data,                         --                 st_sink.data
			st_sink_valid                              => avalon_st_adapter_out_0_valid,                        --                        .valid
			st_sink_ready                              => avalon_st_adapter_out_0_ready,                        --                        .ready
			st_sink_startofpacket                      => avalon_st_adapter_out_0_startofpacket,                --                        .startofpacket
			st_sink_endofpacket                        => avalon_st_adapter_out_0_endofpacket,                  --                        .endofpacket
			st_sink_empty                              => avalon_st_adapter_out_0_empty,                        --                        .empty
			st_sink_error                              => avalon_st_adapter_out_0_error                         --                        .error
		);

	msgdma_tx : component q_sys_msgdma_tx
		port map (
			mm_read_address                            => msgdma_tx_mm_read_address,                            --                 mm_read.address
			mm_read_read                               => msgdma_tx_mm_read_read,                               --                        .read
			mm_read_byteenable                         => msgdma_tx_mm_read_byteenable,                         --                        .byteenable
			mm_read_readdata                           => msgdma_tx_mm_read_readdata,                           --                        .readdata
			mm_read_waitrequest                        => msgdma_tx_mm_read_waitrequest,                        --                        .waitrequest
			mm_read_readdatavalid                      => msgdma_tx_mm_read_readdatavalid,                      --                        .readdatavalid
			descriptor_read_master_address             => msgdma_tx_descriptor_read_master_address,             --  descriptor_read_master.address
			descriptor_read_master_read                => msgdma_tx_descriptor_read_master_read,                --                        .read
			descriptor_read_master_readdata            => msgdma_tx_descriptor_read_master_readdata,            --                        .readdata
			descriptor_read_master_waitrequest         => msgdma_tx_descriptor_read_master_waitrequest,         --                        .waitrequest
			descriptor_read_master_readdatavalid       => msgdma_tx_descriptor_read_master_readdatavalid,       --                        .readdatavalid
			descriptor_write_master_address            => msgdma_tx_descriptor_write_master_address,            -- descriptor_write_master.address
			descriptor_write_master_write              => msgdma_tx_descriptor_write_master_write,              --                        .write
			descriptor_write_master_byteenable         => msgdma_tx_descriptor_write_master_byteenable,         --                        .byteenable
			descriptor_write_master_writedata          => msgdma_tx_descriptor_write_master_writedata,          --                        .writedata
			descriptor_write_master_waitrequest        => msgdma_tx_descriptor_write_master_waitrequest,        --                        .waitrequest
			descriptor_write_master_response           => msgdma_tx_descriptor_write_master_response,           --                        .response
			descriptor_write_master_writeresponsevalid => msgdma_tx_descriptor_write_master_writeresponsevalid, --                        .writeresponsevalid
			clock_clk                                  => sll_hyperbus_controller_top_0_o_av_out_clk_clk,       --                   clock.clk
			reset_n_reset_n                            => sll_hyperbus_controller_top_0_o_av_out_rstn_reset,    --                 reset_n.reset_n
			csr_writedata                              => mm_interconnect_1_msgdma_tx_csr_writedata,            --                     csr.writedata
			csr_write                                  => mm_interconnect_1_msgdma_tx_csr_write,                --                        .write
			csr_byteenable                             => mm_interconnect_1_msgdma_tx_csr_byteenable,           --                        .byteenable
			csr_readdata                               => mm_interconnect_1_msgdma_tx_csr_readdata,             --                        .readdata
			csr_read                                   => mm_interconnect_1_msgdma_tx_csr_read,                 --                        .read
			csr_address                                => mm_interconnect_1_msgdma_tx_csr_address,              --                        .address
			prefetcher_csr_address                     => mm_interconnect_1_msgdma_tx_prefetcher_csr_address,   --          prefetcher_csr.address
			prefetcher_csr_read                        => mm_interconnect_1_msgdma_tx_prefetcher_csr_read,      --                        .read
			prefetcher_csr_write                       => mm_interconnect_1_msgdma_tx_prefetcher_csr_write,     --                        .write
			prefetcher_csr_writedata                   => mm_interconnect_1_msgdma_tx_prefetcher_csr_writedata, --                        .writedata
			prefetcher_csr_readdata                    => mm_interconnect_1_msgdma_tx_prefetcher_csr_readdata,  --                        .readdata
			csr_irq_irq                                => irq_mapper_receiver1_irq,                             --                 csr_irq.irq
			st_source_data                             => msgdma_tx_st_source_data,                             --               st_source.data
			st_source_valid                            => msgdma_tx_st_source_valid,                            --                        .valid
			st_source_ready                            => msgdma_tx_st_source_ready,                            --                        .ready
			st_source_startofpacket                    => msgdma_tx_st_source_startofpacket,                    --                        .startofpacket
			st_source_endofpacket                      => msgdma_tx_st_source_endofpacket,                      --                        .endofpacket
			st_source_empty                            => msgdma_tx_st_source_empty,                            --                        .empty
			st_source_error                            => msgdma_tx_st_source_error                             --                        .error
		);

	onchip_ram : component q_sys_onchip_ram
		port map (
			clk        => sll_hyperbus_controller_top_0_o_av_out_clk_clk, --   clk1.clk
			address    => mm_interconnect_0_onchip_ram_s1_address,        --     s1.address
			clken      => mm_interconnect_0_onchip_ram_s1_clken,          --       .clken
			chipselect => mm_interconnect_0_onchip_ram_s1_chipselect,     --       .chipselect
			write      => mm_interconnect_0_onchip_ram_s1_write,          --       .write
			readdata   => mm_interconnect_0_onchip_ram_s1_readdata,       --       .readdata
			writedata  => mm_interconnect_0_onchip_ram_s1_writedata,      --       .writedata
			byteenable => mm_interconnect_0_onchip_ram_s1_byteenable,     --       .byteenable
			reset      => rst_controller_reset_out_reset,                 -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,             --       .reset_req
			freeze     => '0'                                             -- (terminated)
		);

	opencores_i2c_0 : component opencores_i2c
		generic map (
			FIXED_PRESCALE => 5
		)
		port map (
			wb_clk_i   => sll_hyperbus_controller_top_0_o_av_out_clk_clk,              --            clock.clk
			wb_rst_i   => sll_hyperbus_controller_top_0_o_av_out_rstn_reset_ports_inv, --      clock_reset.reset
			scl_pad_io => opencores_i2c_scl_pad_io,                                    --         export_0.export
			sda_pad_io => opencores_i2c_sda_pad_io,                                    --                 .export
			wb_adr_i   => mm_interconnect_1_opencores_i2c_0_avalon_slave_0_address,    --   avalon_slave_0.address
			wb_dat_i   => mm_interconnect_1_opencores_i2c_0_avalon_slave_0_writedata,  --                 .writedata
			wb_dat_o   => mm_interconnect_1_opencores_i2c_0_avalon_slave_0_readdata,   --                 .readdata
			wb_we_i    => mm_interconnect_1_opencores_i2c_0_avalon_slave_0_write,      --                 .write
			wb_stb_i   => mm_interconnect_1_opencores_i2c_0_avalon_slave_0_chipselect, --                 .chipselect
			wb_ack_o   => opencores_i2c_0_avalon_slave_0_waitrequest,                  --                 .waitrequest_n
			wb_inta_o  => open                                                         -- interrupt_sender.irq
		);

	remote_update : component q_sys_remote_update
		port map (
			avl_csr_write         => mm_interconnect_0_remote_update_avl_csr_write,         -- avl_csr.write
			avl_csr_read          => mm_interconnect_0_remote_update_avl_csr_read,          --        .read
			avl_csr_writedata     => mm_interconnect_0_remote_update_avl_csr_writedata,     --        .writedata
			avl_csr_readdata      => mm_interconnect_0_remote_update_avl_csr_readdata,      --        .readdata
			avl_csr_readdatavalid => mm_interconnect_0_remote_update_avl_csr_readdatavalid, --        .readdatavalid
			avl_csr_waitrequest   => mm_interconnect_0_remote_update_avl_csr_waitrequest,   --        .waitrequest
			avl_csr_address       => mm_interconnect_0_remote_update_avl_csr_address,       --        .address
			clock_clk             => clock_bridge_0_in_clk_clk,                             --   clock.clk
			reset_reset           => rst_controller_002_reset_out_reset                     --   reset.reset
		);

	sll_hyperbus_controller_top_0 : component sll_hyperbus_controller_top
		generic map (
			g_iavs0_addr_width         => 22,
			g_iavs0_data_width         => 32,
			g_iavs0_av_numsymbols      => 4,
			g_iavs0_burstcount_width   => 4,
			g_iavs0_linewrap_burst     => 1,
			g_iavs0_register_rdata     => 0,
			g_iavs0_register_wdata     => 0,
			g_include_reg_avalon       => 0,
			g_include_internal_pll     => 1,
			g_input_clk_freq_in_mhz    => 50,
			g_hyperbus_freq_in_mhz     => 150,
			g_iavs_freq_in_mhz         => 75,
			g_same_iavs_hyperbus_clk   => 0,
			g_config_rd_buffer_as_sram => 1,
			g_config_wr_buffer_as_sram => 1,
			g_device_family            => "Cyclone 10 LP",
			g_num_chipselect           => 2,
			g_dev0_config              => "00000000000000000000000000000000",
			g_dev1_config              => "10001111000111110000000001000001",
			g_dev0_timing              => "00000000000000000000000000000000",
			g_dev1_timing              => "00000000000001100111000100100001",
			g_include_dual_rwds_pin    => 0,
			g_dqin_rdata_width         => 8
		)
		port map (
			in_clk               => hbus_clk_clk,                                                        --        in_clk.clk
			i_ext_rstn           => rst_controller_003_reset_out_reset_ports_inv,                        --    i_ext_rstn.reset_n
			i_iavs0_clk          => sll_hyperbus_controller_top_0_o_av_out_clk_clk,                      --   i_iavs0_clk.clk
			i_iavs0_rstn         => sll_hyperbus_controller_top_0_o_av_out_rstn_reset,                   --  i_iavs0_rstn.reset_n
			i_iavs0_addr         => mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_address,       --         iavs0.address
			i_iavs0_burstcount   => mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_burstcount,    --              .burstcount
			o_iavs0_wait_request => mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_waitrequest,   --              .waitrequest
			i_iavs0_do_wr        => mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_write,         --              .write
			i_iavs0_byteenable   => mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_byteenable,    --              .byteenable
			i_iavs0_wdata        => mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_writedata,     --              .writedata
			i_iavs0_do_rd        => mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_read,          --              .read
			o_iavs0_rdata        => mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_readdata,      --              .readdata
			o_iavs0_rdata_valid  => mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_readdatavalid, --              .readdatavalid
			HB_RSTn              => hyperbus_controller_top_HB_RSTn,                                     --    Conduit_IO.HB_RSTn
			HB_CLK0              => hyperbus_controller_top_HB_CLK0,                                     --              .HB_CLK0
			HB_CLK0n             => hyperbus_controller_top_HB_CLK0n,                                    --              .HB_CLK0n
			HB_CLK1              => hyperbus_controller_top_HB_CLK1,                                     --              .HB_CLK1
			HB_CLK1n             => hyperbus_controller_top_HB_CLK1n,                                    --              .HB_CLK1n
			HB_CS0n              => hyperbus_controller_top_HB_CS0n,                                     --              .HB_CS0n
			HB_CS1n              => hyperbus_controller_top_HB_CS1n,                                     --              .HB_CS1n
			HB_WPn               => hyperbus_controller_top_HB_WPn,                                      --              .HB_WPn
			HB_RWDS              => hyperbus_controller_top_HB_RWDS,                                     --              .HB_RWDS
			HB_dq                => hyperbus_controller_top_HB_dq,                                       --              .HB_dq
			HB_RSTOn             => hyperbus_controller_top_HB_RSTOn,                                    --              .HB_RSTOn
			HB_INTn              => hyperbus_controller_top_HB_INTn,                                     --              .HB_INTn
			o_av_out_clk         => sll_hyperbus_controller_top_0_o_av_out_clk_clk,                      --  o_av_out_clk.clk
			o_av_out_rstn        => sll_hyperbus_controller_top_0_o_av_out_rstn_reset,                   -- o_av_out_rstn.reset_n
			o_iavs0_resp         => open,                                                                --   (terminated)
			i_iavsr_addr         => "000",                                                               --   (terminated)
			i_iavsr_do_wr        => '0',                                                                 --   (terminated)
			i_iavsr_do_rd        => '0',                                                                 --   (terminated)
			i_iavsr_wdata        => "00000000000000000000000000000000",                                  --   (terminated)
			o_iavsr_rdata        => open                                                                 --   (terminated)
		);

	sys_clk_timer : component q_sys_sys_clk_timer
		port map (
			clk        => sll_hyperbus_controller_top_0_o_av_out_clk_clk,     --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,           -- reset.reset_n
			address    => mm_interconnect_1_sys_clk_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_1_sys_clk_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_1_sys_clk_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_1_sys_clk_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_1_sys_clk_timer_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver3_irq                            --   irq.irq
		);

	sysid : component q_sys_sysid
		port map (
			clock    => sll_hyperbus_controller_top_0_o_av_out_clk_clk,   --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,         --         reset.reset_n
			readdata => mm_interconnect_1_sysid_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_1_sysid_control_slave_address(0)  --              .address
		);

	user_dipsw : component q_sys_user_dipsw
		port map (
			clk      => sll_hyperbus_controller_top_0_o_av_out_clk_clk,    --                 clk.clk
			reset_n  => sll_hyperbus_controller_top_0_o_av_out_rstn_reset, --               reset.reset_n
			address  => mm_interconnect_1_user_dipsw_s1_address,           --                  s1.address
			readdata => mm_interconnect_1_user_dipsw_s1_readdata,          --                    .readdata
			in_port  => user_dipsw_external_connection_export              -- external_connection.export
		);

	user_pb : component q_sys_user_dipsw
		port map (
			clk      => sll_hyperbus_controller_top_0_o_av_out_clk_clk,    --                 clk.clk
			reset_n  => sll_hyperbus_controller_top_0_o_av_out_rstn_reset, --               reset.reset_n
			address  => mm_interconnect_1_user_pb_s1_address,              --                  s1.address
			readdata => mm_interconnect_1_user_pb_s1_readdata,             --                    .readdata
			in_port  => user_pb_external_connection_export                 -- external_connection.export
		);

	userhw_0 : component userhw
		port map (
			clk       => sll_hyperbus_controller_top_0_o_av_out_clk_clk,              --          clock.clk
			read      => mm_interconnect_1_userhw_0_avalon_slave_0_read,              -- avalon_slave_0.read
			write     => mm_interconnect_1_userhw_0_avalon_slave_0_write,             --               .write
			address   => mm_interconnect_1_userhw_0_avalon_slave_0_address,           --               .address
			writedata => mm_interconnect_1_userhw_0_avalon_slave_0_writedata,         --               .writedata
			readdata  => mm_interconnect_1_userhw_0_avalon_slave_0_readdata,          --               .readdata
			rst       => sll_hyperbus_controller_top_0_o_av_out_rstn_reset_ports_inv  --     reset_sink.reset
		);

	mm_interconnect_0 : component q_sys_mm_interconnect_0
		port map (
			clock_bridge_0_out_clk_clk                                             => clock_bridge_0_in_clk_clk,                                           --                                           clock_bridge_0_out_clk.clk
			sll_hyperbus_controller_top_0_o_av_out_clk_clk                         => sll_hyperbus_controller_top_0_o_av_out_clk_clk,                      --                       sll_hyperbus_controller_top_0_o_av_out_clk.clk
			cpu_reset_reset_bridge_in_reset_reset                                  => rst_controller_reset_out_reset,                                      --                                  cpu_reset_reset_bridge_in_reset.reset
			ext_epcq_flash_reset_reset_bridge_in_reset_reset                       => rst_controller_002_reset_out_reset,                                  --                       ext_epcq_flash_reset_reset_bridge_in_reset.reset
			sll_hyperbus_controller_top_0_i_iavs0_rstn_reset_bridge_in_reset_reset => sll_hyperbus_controller_top_0_o_av_out_rstn_reset_ports_inv,         -- sll_hyperbus_controller_top_0_i_iavs0_rstn_reset_bridge_in_reset.reset
			cpu_data_master_address                                                => cpu_data_master_address,                                             --                                                  cpu_data_master.address
			cpu_data_master_waitrequest                                            => cpu_data_master_waitrequest,                                         --                                                                 .waitrequest
			cpu_data_master_burstcount                                             => cpu_data_master_burstcount,                                          --                                                                 .burstcount
			cpu_data_master_byteenable                                             => cpu_data_master_byteenable,                                          --                                                                 .byteenable
			cpu_data_master_read                                                   => cpu_data_master_read,                                                --                                                                 .read
			cpu_data_master_readdata                                               => cpu_data_master_readdata,                                            --                                                                 .readdata
			cpu_data_master_readdatavalid                                          => cpu_data_master_readdatavalid,                                       --                                                                 .readdatavalid
			cpu_data_master_write                                                  => cpu_data_master_write,                                               --                                                                 .write
			cpu_data_master_writedata                                              => cpu_data_master_writedata,                                           --                                                                 .writedata
			cpu_data_master_debugaccess                                            => cpu_data_master_debugaccess,                                         --                                                                 .debugaccess
			cpu_instruction_master_address                                         => cpu_instruction_master_address,                                      --                                           cpu_instruction_master.address
			cpu_instruction_master_waitrequest                                     => cpu_instruction_master_waitrequest,                                  --                                                                 .waitrequest
			cpu_instruction_master_burstcount                                      => cpu_instruction_master_burstcount,                                   --                                                                 .burstcount
			cpu_instruction_master_read                                            => cpu_instruction_master_read,                                         --                                                                 .read
			cpu_instruction_master_readdata                                        => cpu_instruction_master_readdata,                                     --                                                                 .readdata
			cpu_instruction_master_readdatavalid                                   => cpu_instruction_master_readdatavalid,                                --                                                                 .readdatavalid
			msgdma_rx_mm_write_address                                             => msgdma_rx_mm_write_address,                                          --                                               msgdma_rx_mm_write.address
			msgdma_rx_mm_write_waitrequest                                         => msgdma_rx_mm_write_waitrequest,                                      --                                                                 .waitrequest
			msgdma_rx_mm_write_byteenable                                          => msgdma_rx_mm_write_byteenable,                                       --                                                                 .byteenable
			msgdma_rx_mm_write_write                                               => msgdma_rx_mm_write_write,                                            --                                                                 .write
			msgdma_rx_mm_write_writedata                                           => msgdma_rx_mm_write_writedata,                                        --                                                                 .writedata
			msgdma_tx_mm_read_address                                              => msgdma_tx_mm_read_address,                                           --                                                msgdma_tx_mm_read.address
			msgdma_tx_mm_read_waitrequest                                          => msgdma_tx_mm_read_waitrequest,                                       --                                                                 .waitrequest
			msgdma_tx_mm_read_byteenable                                           => msgdma_tx_mm_read_byteenable,                                        --                                                                 .byteenable
			msgdma_tx_mm_read_read                                                 => msgdma_tx_mm_read_read,                                              --                                                                 .read
			msgdma_tx_mm_read_readdata                                             => msgdma_tx_mm_read_readdata,                                          --                                                                 .readdata
			msgdma_tx_mm_read_readdatavalid                                        => msgdma_tx_mm_read_readdatavalid,                                     --                                                                 .readdatavalid
			cpu_debug_mem_slave_address                                            => mm_interconnect_0_cpu_debug_mem_slave_address,                       --                                              cpu_debug_mem_slave.address
			cpu_debug_mem_slave_write                                              => mm_interconnect_0_cpu_debug_mem_slave_write,                         --                                                                 .write
			cpu_debug_mem_slave_read                                               => mm_interconnect_0_cpu_debug_mem_slave_read,                          --                                                                 .read
			cpu_debug_mem_slave_readdata                                           => mm_interconnect_0_cpu_debug_mem_slave_readdata,                      --                                                                 .readdata
			cpu_debug_mem_slave_writedata                                          => mm_interconnect_0_cpu_debug_mem_slave_writedata,                     --                                                                 .writedata
			cpu_debug_mem_slave_byteenable                                         => mm_interconnect_0_cpu_debug_mem_slave_byteenable,                    --                                                                 .byteenable
			cpu_debug_mem_slave_waitrequest                                        => mm_interconnect_0_cpu_debug_mem_slave_waitrequest,                   --                                                                 .waitrequest
			cpu_debug_mem_slave_debugaccess                                        => mm_interconnect_0_cpu_debug_mem_slave_debugaccess,                   --                                                                 .debugaccess
			ext_epcq_flash_avl_csr_address                                         => mm_interconnect_0_ext_epcq_flash_avl_csr_address,                    --                                           ext_epcq_flash_avl_csr.address
			ext_epcq_flash_avl_csr_write                                           => mm_interconnect_0_ext_epcq_flash_avl_csr_write,                      --                                                                 .write
			ext_epcq_flash_avl_csr_read                                            => mm_interconnect_0_ext_epcq_flash_avl_csr_read,                       --                                                                 .read
			ext_epcq_flash_avl_csr_readdata                                        => mm_interconnect_0_ext_epcq_flash_avl_csr_readdata,                   --                                                                 .readdata
			ext_epcq_flash_avl_csr_writedata                                       => mm_interconnect_0_ext_epcq_flash_avl_csr_writedata,                  --                                                                 .writedata
			ext_epcq_flash_avl_csr_readdatavalid                                   => mm_interconnect_0_ext_epcq_flash_avl_csr_readdatavalid,              --                                                                 .readdatavalid
			ext_epcq_flash_avl_csr_waitrequest                                     => mm_interconnect_0_ext_epcq_flash_avl_csr_waitrequest,                --                                                                 .waitrequest
			ext_epcq_flash_avl_mem_address                                         => mm_interconnect_0_ext_epcq_flash_avl_mem_address,                    --                                           ext_epcq_flash_avl_mem.address
			ext_epcq_flash_avl_mem_write                                           => mm_interconnect_0_ext_epcq_flash_avl_mem_write,                      --                                                                 .write
			ext_epcq_flash_avl_mem_read                                            => mm_interconnect_0_ext_epcq_flash_avl_mem_read,                       --                                                                 .read
			ext_epcq_flash_avl_mem_readdata                                        => mm_interconnect_0_ext_epcq_flash_avl_mem_readdata,                   --                                                                 .readdata
			ext_epcq_flash_avl_mem_writedata                                       => mm_interconnect_0_ext_epcq_flash_avl_mem_writedata,                  --                                                                 .writedata
			ext_epcq_flash_avl_mem_burstcount                                      => mm_interconnect_0_ext_epcq_flash_avl_mem_burstcount,                 --                                                                 .burstcount
			ext_epcq_flash_avl_mem_byteenable                                      => mm_interconnect_0_ext_epcq_flash_avl_mem_byteenable,                 --                                                                 .byteenable
			ext_epcq_flash_avl_mem_readdatavalid                                   => mm_interconnect_0_ext_epcq_flash_avl_mem_readdatavalid,              --                                                                 .readdatavalid
			ext_epcq_flash_avl_mem_waitrequest                                     => mm_interconnect_0_ext_epcq_flash_avl_mem_waitrequest,                --                                                                 .waitrequest
			mm_bridge_0_s0_address                                                 => mm_interconnect_0_mm_bridge_0_s0_address,                            --                                                   mm_bridge_0_s0.address
			mm_bridge_0_s0_write                                                   => mm_interconnect_0_mm_bridge_0_s0_write,                              --                                                                 .write
			mm_bridge_0_s0_read                                                    => mm_interconnect_0_mm_bridge_0_s0_read,                               --                                                                 .read
			mm_bridge_0_s0_readdata                                                => mm_interconnect_0_mm_bridge_0_s0_readdata,                           --                                                                 .readdata
			mm_bridge_0_s0_writedata                                               => mm_interconnect_0_mm_bridge_0_s0_writedata,                          --                                                                 .writedata
			mm_bridge_0_s0_burstcount                                              => mm_interconnect_0_mm_bridge_0_s0_burstcount,                         --                                                                 .burstcount
			mm_bridge_0_s0_byteenable                                              => mm_interconnect_0_mm_bridge_0_s0_byteenable,                         --                                                                 .byteenable
			mm_bridge_0_s0_readdatavalid                                           => mm_interconnect_0_mm_bridge_0_s0_readdatavalid,                      --                                                                 .readdatavalid
			mm_bridge_0_s0_waitrequest                                             => mm_interconnect_0_mm_bridge_0_s0_waitrequest,                        --                                                                 .waitrequest
			mm_bridge_0_s0_debugaccess                                             => mm_interconnect_0_mm_bridge_0_s0_debugaccess,                        --                                                                 .debugaccess
			onchip_ram_s1_address                                                  => mm_interconnect_0_onchip_ram_s1_address,                             --                                                    onchip_ram_s1.address
			onchip_ram_s1_write                                                    => mm_interconnect_0_onchip_ram_s1_write,                               --                                                                 .write
			onchip_ram_s1_readdata                                                 => mm_interconnect_0_onchip_ram_s1_readdata,                            --                                                                 .readdata
			onchip_ram_s1_writedata                                                => mm_interconnect_0_onchip_ram_s1_writedata,                           --                                                                 .writedata
			onchip_ram_s1_byteenable                                               => mm_interconnect_0_onchip_ram_s1_byteenable,                          --                                                                 .byteenable
			onchip_ram_s1_chipselect                                               => mm_interconnect_0_onchip_ram_s1_chipselect,                          --                                                                 .chipselect
			onchip_ram_s1_clken                                                    => mm_interconnect_0_onchip_ram_s1_clken,                               --                                                                 .clken
			remote_update_avl_csr_address                                          => mm_interconnect_0_remote_update_avl_csr_address,                     --                                            remote_update_avl_csr.address
			remote_update_avl_csr_write                                            => mm_interconnect_0_remote_update_avl_csr_write,                       --                                                                 .write
			remote_update_avl_csr_read                                             => mm_interconnect_0_remote_update_avl_csr_read,                        --                                                                 .read
			remote_update_avl_csr_readdata                                         => mm_interconnect_0_remote_update_avl_csr_readdata,                    --                                                                 .readdata
			remote_update_avl_csr_writedata                                        => mm_interconnect_0_remote_update_avl_csr_writedata,                   --                                                                 .writedata
			remote_update_avl_csr_readdatavalid                                    => mm_interconnect_0_remote_update_avl_csr_readdatavalid,               --                                                                 .readdatavalid
			remote_update_avl_csr_waitrequest                                      => mm_interconnect_0_remote_update_avl_csr_waitrequest,                 --                                                                 .waitrequest
			sll_hyperbus_controller_top_0_iavs0_address                            => mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_address,       --                              sll_hyperbus_controller_top_0_iavs0.address
			sll_hyperbus_controller_top_0_iavs0_write                              => mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_write,         --                                                                 .write
			sll_hyperbus_controller_top_0_iavs0_read                               => mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_read,          --                                                                 .read
			sll_hyperbus_controller_top_0_iavs0_readdata                           => mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_readdata,      --                                                                 .readdata
			sll_hyperbus_controller_top_0_iavs0_writedata                          => mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_writedata,     --                                                                 .writedata
			sll_hyperbus_controller_top_0_iavs0_burstcount                         => mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_burstcount,    --                                                                 .burstcount
			sll_hyperbus_controller_top_0_iavs0_byteenable                         => mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_byteenable,    --                                                                 .byteenable
			sll_hyperbus_controller_top_0_iavs0_readdatavalid                      => mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_readdatavalid, --                                                                 .readdatavalid
			sll_hyperbus_controller_top_0_iavs0_waitrequest                        => mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_waitrequest    --                                                                 .waitrequest
		);

	mm_interconnect_1 : component q_sys_mm_interconnect_1
		port map (
			sll_hyperbus_controller_top_0_o_av_out_clk_clk       => sll_hyperbus_controller_top_0_o_av_out_clk_clk,              --     sll_hyperbus_controller_top_0_o_av_out_clk.clk
			descriptor_memory_reset1_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                              -- descriptor_memory_reset1_reset_bridge_in_reset.reset
			msgdma_rx_reset_n_reset_bridge_in_reset_reset        => sll_hyperbus_controller_top_0_o_av_out_rstn_reset_ports_inv, --        msgdma_rx_reset_n_reset_bridge_in_reset.reset
			mm_bridge_0_m0_address                               => mm_bridge_0_m0_address,                                      --                                 mm_bridge_0_m0.address
			mm_bridge_0_m0_waitrequest                           => mm_bridge_0_m0_waitrequest,                                  --                                               .waitrequest
			mm_bridge_0_m0_burstcount                            => mm_bridge_0_m0_burstcount,                                   --                                               .burstcount
			mm_bridge_0_m0_byteenable                            => mm_bridge_0_m0_byteenable,                                   --                                               .byteenable
			mm_bridge_0_m0_read                                  => mm_bridge_0_m0_read,                                         --                                               .read
			mm_bridge_0_m0_readdata                              => mm_bridge_0_m0_readdata,                                     --                                               .readdata
			mm_bridge_0_m0_readdatavalid                         => mm_bridge_0_m0_readdatavalid,                                --                                               .readdatavalid
			mm_bridge_0_m0_write                                 => mm_bridge_0_m0_write,                                        --                                               .write
			mm_bridge_0_m0_writedata                             => mm_bridge_0_m0_writedata,                                    --                                               .writedata
			mm_bridge_0_m0_debugaccess                           => mm_bridge_0_m0_debugaccess,                                  --                                               .debugaccess
			msgdma_rx_descriptor_read_master_address             => msgdma_rx_descriptor_read_master_address,                    --               msgdma_rx_descriptor_read_master.address
			msgdma_rx_descriptor_read_master_waitrequest         => msgdma_rx_descriptor_read_master_waitrequest,                --                                               .waitrequest
			msgdma_rx_descriptor_read_master_read                => msgdma_rx_descriptor_read_master_read,                       --                                               .read
			msgdma_rx_descriptor_read_master_readdata            => msgdma_rx_descriptor_read_master_readdata,                   --                                               .readdata
			msgdma_rx_descriptor_read_master_readdatavalid       => msgdma_rx_descriptor_read_master_readdatavalid,              --                                               .readdatavalid
			msgdma_rx_descriptor_write_master_address            => msgdma_rx_descriptor_write_master_address,                   --              msgdma_rx_descriptor_write_master.address
			msgdma_rx_descriptor_write_master_waitrequest        => msgdma_rx_descriptor_write_master_waitrequest,               --                                               .waitrequest
			msgdma_rx_descriptor_write_master_byteenable         => msgdma_rx_descriptor_write_master_byteenable,                --                                               .byteenable
			msgdma_rx_descriptor_write_master_write              => msgdma_rx_descriptor_write_master_write,                     --                                               .write
			msgdma_rx_descriptor_write_master_writedata          => msgdma_rx_descriptor_write_master_writedata,                 --                                               .writedata
			msgdma_rx_descriptor_write_master_response           => msgdma_rx_descriptor_write_master_response,                  --                                               .response
			msgdma_rx_descriptor_write_master_writeresponsevalid => msgdma_rx_descriptor_write_master_writeresponsevalid,        --                                               .writeresponsevalid
			msgdma_tx_descriptor_read_master_address             => msgdma_tx_descriptor_read_master_address,                    --               msgdma_tx_descriptor_read_master.address
			msgdma_tx_descriptor_read_master_waitrequest         => msgdma_tx_descriptor_read_master_waitrequest,                --                                               .waitrequest
			msgdma_tx_descriptor_read_master_read                => msgdma_tx_descriptor_read_master_read,                       --                                               .read
			msgdma_tx_descriptor_read_master_readdata            => msgdma_tx_descriptor_read_master_readdata,                   --                                               .readdata
			msgdma_tx_descriptor_read_master_readdatavalid       => msgdma_tx_descriptor_read_master_readdatavalid,              --                                               .readdatavalid
			msgdma_tx_descriptor_write_master_address            => msgdma_tx_descriptor_write_master_address,                   --              msgdma_tx_descriptor_write_master.address
			msgdma_tx_descriptor_write_master_waitrequest        => msgdma_tx_descriptor_write_master_waitrequest,               --                                               .waitrequest
			msgdma_tx_descriptor_write_master_byteenable         => msgdma_tx_descriptor_write_master_byteenable,                --                                               .byteenable
			msgdma_tx_descriptor_write_master_write              => msgdma_tx_descriptor_write_master_write,                     --                                               .write
			msgdma_tx_descriptor_write_master_writedata          => msgdma_tx_descriptor_write_master_writedata,                 --                                               .writedata
			msgdma_tx_descriptor_write_master_response           => msgdma_tx_descriptor_write_master_response,                  --                                               .response
			msgdma_tx_descriptor_write_master_writeresponsevalid => msgdma_tx_descriptor_write_master_writeresponsevalid,        --                                               .writeresponsevalid
			descriptor_memory_s1_address                         => mm_interconnect_1_descriptor_memory_s1_address,              --                           descriptor_memory_s1.address
			descriptor_memory_s1_write                           => mm_interconnect_1_descriptor_memory_s1_write,                --                                               .write
			descriptor_memory_s1_readdata                        => mm_interconnect_1_descriptor_memory_s1_readdata,             --                                               .readdata
			descriptor_memory_s1_writedata                       => mm_interconnect_1_descriptor_memory_s1_writedata,            --                                               .writedata
			descriptor_memory_s1_byteenable                      => mm_interconnect_1_descriptor_memory_s1_byteenable,           --                                               .byteenable
			descriptor_memory_s1_chipselect                      => mm_interconnect_1_descriptor_memory_s1_chipselect,           --                                               .chipselect
			descriptor_memory_s1_clken                           => mm_interconnect_1_descriptor_memory_s1_clken,                --                                               .clken
			eth_tse_control_port_address                         => mm_interconnect_1_eth_tse_control_port_address,              --                           eth_tse_control_port.address
			eth_tse_control_port_write                           => mm_interconnect_1_eth_tse_control_port_write,                --                                               .write
			eth_tse_control_port_read                            => mm_interconnect_1_eth_tse_control_port_read,                 --                                               .read
			eth_tse_control_port_readdata                        => mm_interconnect_1_eth_tse_control_port_readdata,             --                                               .readdata
			eth_tse_control_port_writedata                       => mm_interconnect_1_eth_tse_control_port_writedata,            --                                               .writedata
			eth_tse_control_port_waitrequest                     => mm_interconnect_1_eth_tse_control_port_waitrequest,          --                                               .waitrequest
			jtag_uart_avalon_jtag_slave_address                  => mm_interconnect_1_jtag_uart_avalon_jtag_slave_address,       --                    jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write                    => mm_interconnect_1_jtag_uart_avalon_jtag_slave_write,         --                                               .write
			jtag_uart_avalon_jtag_slave_read                     => mm_interconnect_1_jtag_uart_avalon_jtag_slave_read,          --                                               .read
			jtag_uart_avalon_jtag_slave_readdata                 => mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata,      --                                               .readdata
			jtag_uart_avalon_jtag_slave_writedata                => mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata,     --                                               .writedata
			jtag_uart_avalon_jtag_slave_waitrequest              => mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest,   --                                               .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect               => mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect,    --                                               .chipselect
			led_pio_s1_address                                   => mm_interconnect_1_led_pio_s1_address,                        --                                     led_pio_s1.address
			led_pio_s1_write                                     => mm_interconnect_1_led_pio_s1_write,                          --                                               .write
			led_pio_s1_readdata                                  => mm_interconnect_1_led_pio_s1_readdata,                       --                                               .readdata
			led_pio_s1_writedata                                 => mm_interconnect_1_led_pio_s1_writedata,                      --                                               .writedata
			led_pio_s1_chipselect                                => mm_interconnect_1_led_pio_s1_chipselect,                     --                                               .chipselect
			msgdma_rx_csr_address                                => mm_interconnect_1_msgdma_rx_csr_address,                     --                                  msgdma_rx_csr.address
			msgdma_rx_csr_write                                  => mm_interconnect_1_msgdma_rx_csr_write,                       --                                               .write
			msgdma_rx_csr_read                                   => mm_interconnect_1_msgdma_rx_csr_read,                        --                                               .read
			msgdma_rx_csr_readdata                               => mm_interconnect_1_msgdma_rx_csr_readdata,                    --                                               .readdata
			msgdma_rx_csr_writedata                              => mm_interconnect_1_msgdma_rx_csr_writedata,                   --                                               .writedata
			msgdma_rx_csr_byteenable                             => mm_interconnect_1_msgdma_rx_csr_byteenable,                  --                                               .byteenable
			msgdma_rx_prefetcher_csr_address                     => mm_interconnect_1_msgdma_rx_prefetcher_csr_address,          --                       msgdma_rx_prefetcher_csr.address
			msgdma_rx_prefetcher_csr_write                       => mm_interconnect_1_msgdma_rx_prefetcher_csr_write,            --                                               .write
			msgdma_rx_prefetcher_csr_read                        => mm_interconnect_1_msgdma_rx_prefetcher_csr_read,             --                                               .read
			msgdma_rx_prefetcher_csr_readdata                    => mm_interconnect_1_msgdma_rx_prefetcher_csr_readdata,         --                                               .readdata
			msgdma_rx_prefetcher_csr_writedata                   => mm_interconnect_1_msgdma_rx_prefetcher_csr_writedata,        --                                               .writedata
			msgdma_tx_csr_address                                => mm_interconnect_1_msgdma_tx_csr_address,                     --                                  msgdma_tx_csr.address
			msgdma_tx_csr_write                                  => mm_interconnect_1_msgdma_tx_csr_write,                       --                                               .write
			msgdma_tx_csr_read                                   => mm_interconnect_1_msgdma_tx_csr_read,                        --                                               .read
			msgdma_tx_csr_readdata                               => mm_interconnect_1_msgdma_tx_csr_readdata,                    --                                               .readdata
			msgdma_tx_csr_writedata                              => mm_interconnect_1_msgdma_tx_csr_writedata,                   --                                               .writedata
			msgdma_tx_csr_byteenable                             => mm_interconnect_1_msgdma_tx_csr_byteenable,                  --                                               .byteenable
			msgdma_tx_prefetcher_csr_address                     => mm_interconnect_1_msgdma_tx_prefetcher_csr_address,          --                       msgdma_tx_prefetcher_csr.address
			msgdma_tx_prefetcher_csr_write                       => mm_interconnect_1_msgdma_tx_prefetcher_csr_write,            --                                               .write
			msgdma_tx_prefetcher_csr_read                        => mm_interconnect_1_msgdma_tx_prefetcher_csr_read,             --                                               .read
			msgdma_tx_prefetcher_csr_readdata                    => mm_interconnect_1_msgdma_tx_prefetcher_csr_readdata,         --                                               .readdata
			msgdma_tx_prefetcher_csr_writedata                   => mm_interconnect_1_msgdma_tx_prefetcher_csr_writedata,        --                                               .writedata
			opencores_i2c_0_avalon_slave_0_address               => mm_interconnect_1_opencores_i2c_0_avalon_slave_0_address,    --                 opencores_i2c_0_avalon_slave_0.address
			opencores_i2c_0_avalon_slave_0_write                 => mm_interconnect_1_opencores_i2c_0_avalon_slave_0_write,      --                                               .write
			opencores_i2c_0_avalon_slave_0_readdata              => mm_interconnect_1_opencores_i2c_0_avalon_slave_0_readdata,   --                                               .readdata
			opencores_i2c_0_avalon_slave_0_writedata             => mm_interconnect_1_opencores_i2c_0_avalon_slave_0_writedata,  --                                               .writedata
			opencores_i2c_0_avalon_slave_0_waitrequest           => mm_interconnect_1_opencores_i2c_0_avalon_slave_0_inv,        --                                               .waitrequest
			opencores_i2c_0_avalon_slave_0_chipselect            => mm_interconnect_1_opencores_i2c_0_avalon_slave_0_chipselect, --                                               .chipselect
			sys_clk_timer_s1_address                             => mm_interconnect_1_sys_clk_timer_s1_address,                  --                               sys_clk_timer_s1.address
			sys_clk_timer_s1_write                               => mm_interconnect_1_sys_clk_timer_s1_write,                    --                                               .write
			sys_clk_timer_s1_readdata                            => mm_interconnect_1_sys_clk_timer_s1_readdata,                 --                                               .readdata
			sys_clk_timer_s1_writedata                           => mm_interconnect_1_sys_clk_timer_s1_writedata,                --                                               .writedata
			sys_clk_timer_s1_chipselect                          => mm_interconnect_1_sys_clk_timer_s1_chipselect,               --                                               .chipselect
			sysid_control_slave_address                          => mm_interconnect_1_sysid_control_slave_address,               --                            sysid_control_slave.address
			sysid_control_slave_readdata                         => mm_interconnect_1_sysid_control_slave_readdata,              --                                               .readdata
			user_dipsw_s1_address                                => mm_interconnect_1_user_dipsw_s1_address,                     --                                  user_dipsw_s1.address
			user_dipsw_s1_readdata                               => mm_interconnect_1_user_dipsw_s1_readdata,                    --                                               .readdata
			user_pb_s1_address                                   => mm_interconnect_1_user_pb_s1_address,                        --                                     user_pb_s1.address
			user_pb_s1_readdata                                  => mm_interconnect_1_user_pb_s1_readdata,                       --                                               .readdata
			userhw_0_avalon_slave_0_address                      => mm_interconnect_1_userhw_0_avalon_slave_0_address,           --                        userhw_0_avalon_slave_0.address
			userhw_0_avalon_slave_0_write                        => mm_interconnect_1_userhw_0_avalon_slave_0_write,             --                                               .write
			userhw_0_avalon_slave_0_read                         => mm_interconnect_1_userhw_0_avalon_slave_0_read,              --                                               .read
			userhw_0_avalon_slave_0_readdata                     => mm_interconnect_1_userhw_0_avalon_slave_0_readdata,          --                                               .readdata
			userhw_0_avalon_slave_0_writedata                    => mm_interconnect_1_userhw_0_avalon_slave_0_writedata          --                                               .writedata
		);

	irq_mapper : component q_sys_irq_mapper
		port map (
			clk           => sll_hyperbus_controller_top_0_o_av_out_clk_clk, --       clk.clk
			reset         => rst_controller_reset_out_reset,                 -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,                       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,                       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,                       -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,                       -- receiver3.irq
			sender_irq    => cpu_irq_irq                                     --    sender.irq
		);

	avalon_st_adapter : component q_sys_avalon_st_adapter
		generic map (
			inBitsPerSymbol => 8,
			inUsePackets    => 1,
			inDataWidth     => 32,
			inChannelWidth  => 0,
			inErrorWidth    => 6,
			inUseEmptyPort  => 1,
			inUseValid      => 1,
			inUseReady      => 1,
			inReadyLatency  => 2,
			outDataWidth    => 32,
			outChannelWidth => 0,
			outErrorWidth   => 6,
			outUseEmptyPort => 1,
			outUseValid     => 1,
			outUseReady     => 1,
			outReadyLatency => 0
		)
		port map (
			in_clk_0_clk        => sll_hyperbus_controller_top_0_o_av_out_clk_clk, -- in_clk_0.clk
			in_rst_0_reset      => rst_controller_reset_out_reset,                 -- in_rst_0.reset
			in_0_data           => eth_tse_receive_data,                           --     in_0.data
			in_0_valid          => eth_tse_receive_valid,                          --         .valid
			in_0_ready          => eth_tse_receive_ready,                          --         .ready
			in_0_startofpacket  => eth_tse_receive_startofpacket,                  --         .startofpacket
			in_0_endofpacket    => eth_tse_receive_endofpacket,                    --         .endofpacket
			in_0_empty          => eth_tse_receive_empty,                          --         .empty
			in_0_error          => eth_tse_receive_error,                          --         .error
			out_0_data          => avalon_st_adapter_out_0_data,                   --    out_0.data
			out_0_valid         => avalon_st_adapter_out_0_valid,                  --         .valid
			out_0_ready         => avalon_st_adapter_out_0_ready,                  --         .ready
			out_0_startofpacket => avalon_st_adapter_out_0_startofpacket,          --         .startofpacket
			out_0_endofpacket   => avalon_st_adapter_out_0_endofpacket,            --         .endofpacket
			out_0_empty         => avalon_st_adapter_out_0_empty,                  --         .empty
			out_0_error         => avalon_st_adapter_out_0_error                   --         .error
		);

	rst_controller : component q_sys_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => cpu_debug_reset_request_reset,                               -- reset_in0.reset
			reset_in1      => sll_hyperbus_controller_top_0_o_av_out_rstn_reset_ports_inv, -- reset_in1.reset
			clk            => sll_hyperbus_controller_top_0_o_av_out_clk_clk,              --       clk.clk
			reset_out      => rst_controller_reset_out_reset,                              -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,                          --          .reset_req
			reset_req_in0  => '0',                                                         -- (terminated)
			reset_req_in1  => '0',                                                         -- (terminated)
			reset_in2      => '0',                                                         -- (terminated)
			reset_req_in2  => '0',                                                         -- (terminated)
			reset_in3      => '0',                                                         -- (terminated)
			reset_req_in3  => '0',                                                         -- (terminated)
			reset_in4      => '0',                                                         -- (terminated)
			reset_req_in4  => '0',                                                         -- (terminated)
			reset_in5      => '0',                                                         -- (terminated)
			reset_req_in5  => '0',                                                         -- (terminated)
			reset_in6      => '0',                                                         -- (terminated)
			reset_req_in6  => '0',                                                         -- (terminated)
			reset_in7      => '0',                                                         -- (terminated)
			reset_req_in7  => '0',                                                         -- (terminated)
			reset_in8      => '0',                                                         -- (terminated)
			reset_req_in8  => '0',                                                         -- (terminated)
			reset_in9      => '0',                                                         -- (terminated)
			reset_req_in9  => '0',                                                         -- (terminated)
			reset_in10     => '0',                                                         -- (terminated)
			reset_req_in10 => '0',                                                         -- (terminated)
			reset_in11     => '0',                                                         -- (terminated)
			reset_req_in11 => '0',                                                         -- (terminated)
			reset_in12     => '0',                                                         -- (terminated)
			reset_req_in12 => '0',                                                         -- (terminated)
			reset_in13     => '0',                                                         -- (terminated)
			reset_req_in13 => '0',                                                         -- (terminated)
			reset_in14     => '0',                                                         -- (terminated)
			reset_req_in14 => '0',                                                         -- (terminated)
			reset_in15     => '0',                                                         -- (terminated)
			reset_req_in15 => '0'                                                          -- (terminated)
		);

	rst_controller_001 : component q_sys_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_enet_reset_n_ports_inv,       -- reset_in0.reset
			clk            => enet_clk_125m_in_clk,               --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_002 : component q_sys_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => hbus_reset_reset_n_ports_inv,       -- reset_in0.reset
			clk            => clock_bridge_0_in_clk_clk,          --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_003 : component q_sys_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => hbus_reset_reset_n_ports_inv,       -- reset_in0.reset
			clk            => hbus_clk_clk,                       --       clk.clk
			reset_out      => rst_controller_003_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	hbus_reset_reset_n_ports_inv <= not hbus_reset_reset_n;

	reset_enet_reset_n_ports_inv <= not reset_enet_reset_n;

	sll_hyperbus_controller_top_0_o_av_out_rstn_reset_ports_inv <= not sll_hyperbus_controller_top_0_o_av_out_rstn_reset;

	mm_interconnect_1_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_1_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_1_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_1_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_1_opencores_i2c_0_avalon_slave_0_inv <= not opencores_i2c_0_avalon_slave_0_waitrequest;

	mm_interconnect_1_sys_clk_timer_s1_write_ports_inv <= not mm_interconnect_1_sys_clk_timer_s1_write;

	mm_interconnect_1_led_pio_s1_write_ports_inv <= not mm_interconnect_1_led_pio_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_002_reset_out_reset_ports_inv <= not rst_controller_002_reset_out_reset;

	rst_controller_003_reset_out_reset_ports_inv <= not rst_controller_003_reset_out_reset;

end architecture rtl; -- of q_sys
