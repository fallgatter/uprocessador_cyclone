// q_sys.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module q_sys (
		input  wire       clock_bridge_0_in_clk_clk,               //               clock_bridge_0_in_clk.clk
		input  wire       enet_clk_125m_in_clk,                    //                    enet_clk_125m_in.clk
		input  wire       enet_pll_areset_conduit_export,          //             enet_pll_areset_conduit.export
		output wire       enet_pll_c0_125m_clk,                    //                    enet_pll_c0_125m.clk
		output wire       enet_pll_c1_25m_clk,                     //                     enet_pll_c1_25m.clk
		output wire       enet_pll_c2_2m5_clk,                     //                     enet_pll_c2_2m5.clk
		output wire       enet_pll_c3_125m_shift_clk,              //              enet_pll_c3_125m_shift.clk
		output wire       enet_pll_c4_25m_shift_clk,               //               enet_pll_c4_25m_shift.clk
		output wire       enet_pll_locked_conduit_export,          //             enet_pll_locked_conduit.export
		output wire       eth_tse_mac_mdio_connection_mdc,         //         eth_tse_mac_mdio_connection.mdc
		input  wire       eth_tse_mac_mdio_connection_mdio_in,     //                                    .mdio_in
		output wire       eth_tse_mac_mdio_connection_mdio_out,    //                                    .mdio_out
		output wire       eth_tse_mac_mdio_connection_mdio_oen,    //                                    .mdio_oen
		input  wire [3:0] eth_tse_mac_rgmii_connection_rgmii_in,   //        eth_tse_mac_rgmii_connection.rgmii_in
		output wire [3:0] eth_tse_mac_rgmii_connection_rgmii_out,  //                                    .rgmii_out
		input  wire       eth_tse_mac_rgmii_connection_rx_control, //                                    .rx_control
		output wire       eth_tse_mac_rgmii_connection_tx_control, //                                    .tx_control
		input  wire       eth_tse_mac_status_connection_set_10,    //       eth_tse_mac_status_connection.set_10
		input  wire       eth_tse_mac_status_connection_set_1000,  //                                    .set_1000
		output wire       eth_tse_mac_status_connection_eth_mode,  //                                    .eth_mode
		output wire       eth_tse_mac_status_connection_ena_10,    //                                    .ena_10
		input  wire       eth_tse_pcs_mac_rx_clock_connection_clk, // eth_tse_pcs_mac_rx_clock_connection.clk
		input  wire       eth_tse_pcs_mac_tx_clock_connection_clk, // eth_tse_pcs_mac_tx_clock_connection.clk
		input  wire       hbus_clk_clk,                            //                            hbus_clk.clk
		input  wire       hbus_reset_reset_n,                      //                          hbus_reset.reset_n
		output wire       hyperbus_controller_top_HB_RSTn,         //             hyperbus_controller_top.HB_RSTn
		output wire       hyperbus_controller_top_HB_CLK0,         //                                    .HB_CLK0
		output wire       hyperbus_controller_top_HB_CLK0n,        //                                    .HB_CLK0n
		output wire       hyperbus_controller_top_HB_CLK1,         //                                    .HB_CLK1
		output wire       hyperbus_controller_top_HB_CLK1n,        //                                    .HB_CLK1n
		output wire       hyperbus_controller_top_HB_CS0n,         //                                    .HB_CS0n
		output wire       hyperbus_controller_top_HB_CS1n,         //                                    .HB_CS1n
		output wire       hyperbus_controller_top_HB_WPn,          //                                    .HB_WPn
		inout  wire       hyperbus_controller_top_HB_RWDS,         //                                    .HB_RWDS
		inout  wire [7:0] hyperbus_controller_top_HB_dq,           //                                    .HB_dq
		input  wire       hyperbus_controller_top_HB_RSTOn,        //                                    .HB_RSTOn
		input  wire       hyperbus_controller_top_HB_INTn,         //                                    .HB_INTn
		output wire [3:0] led_pio_external_connection_export,      //         led_pio_external_connection.export
		inout  wire       opencores_i2c_scl_pad_io,                //                       opencores_i2c.scl_pad_io
		inout  wire       opencores_i2c_sda_pad_io,                //                                    .sda_pad_io
		input  wire       reset_enet_reset_n,                      //                          reset_enet.reset_n
		input  wire [3:0] user_dipsw_external_connection_export,   //      user_dipsw_external_connection.export
		input  wire [3:0] user_pb_external_connection_export       //         user_pb_external_connection.export
	);

	wire         msgdma_tx_st_source_valid;                                           // msgdma_tx:st_source_valid -> eth_tse:ff_tx_wren
	wire  [31:0] msgdma_tx_st_source_data;                                            // msgdma_tx:st_source_data -> eth_tse:ff_tx_data
	wire         msgdma_tx_st_source_ready;                                           // eth_tse:ff_tx_rdy -> msgdma_tx:st_source_ready
	wire         msgdma_tx_st_source_startofpacket;                                   // msgdma_tx:st_source_startofpacket -> eth_tse:ff_tx_sop
	wire         msgdma_tx_st_source_endofpacket;                                     // msgdma_tx:st_source_endofpacket -> eth_tse:ff_tx_eop
	wire         msgdma_tx_st_source_error;                                           // msgdma_tx:st_source_error -> eth_tse:ff_tx_err
	wire   [1:0] msgdma_tx_st_source_empty;                                           // msgdma_tx:st_source_empty -> eth_tse:ff_tx_mod
	wire         sll_hyperbus_controller_top_0_o_av_out_clk_clk;                      // sll_hyperbus_controller_top_0:o_av_out_clk -> [avalon_st_adapter:in_clk_0_clk, cpu:clk, descriptor_memory:clk, eth_tse:clk, eth_tse:ff_rx_clk, eth_tse:ff_tx_clk, irq_mapper:clk, jtag_uart:clk, led_pio:clk, mm_bridge_0:clk, mm_interconnect_0:sll_hyperbus_controller_top_0_o_av_out_clk_clk, mm_interconnect_1:sll_hyperbus_controller_top_0_o_av_out_clk_clk, msgdma_rx:clock_clk, msgdma_tx:clock_clk, onchip_ram:clk, opencores_i2c_0:wb_clk_i, rst_controller:clk, sll_hyperbus_controller_top_0:i_iavs0_clk, sys_clk_timer:clk, sysid:clock, user_dipsw:clk, user_pb:clk]
	wire         sll_hyperbus_controller_top_0_o_av_out_rstn_reset;                   // sll_hyperbus_controller_top_0:o_av_out_rstn -> [mm_bridge_0:reset, mm_interconnect_0:sll_hyperbus_controller_top_0_i_iavs0_rstn_reset_bridge_in_reset_reset, mm_interconnect_1:msgdma_rx_reset_n_reset_bridge_in_reset_reset, msgdma_rx:reset_n_reset_n, msgdma_tx:reset_n_reset_n, opencores_i2c_0:wb_rst_i, rst_controller:reset_in1, sll_hyperbus_controller_top_0:i_iavs0_rstn, user_dipsw:reset_n, user_pb:reset_n]
	wire  [31:0] cpu_data_master_readdata;                                            // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                                         // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                                         // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [26:0] cpu_data_master_address;                                             // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                          // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                                // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_readdatavalid;                                       // mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	wire         cpu_data_master_write;                                               // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                           // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire   [3:0] cpu_data_master_burstcount;                                          // cpu:d_burstcount -> mm_interconnect_0:cpu_data_master_burstcount
	wire  [31:0] cpu_instruction_master_readdata;                                     // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                                  // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [26:0] cpu_instruction_master_address;                                      // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                         // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         cpu_instruction_master_readdatavalid;                                // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire   [3:0] cpu_instruction_master_burstcount;                                   // cpu:i_burstcount -> mm_interconnect_0:cpu_instruction_master_burstcount
	wire  [31:0] msgdma_tx_mm_read_readdata;                                          // mm_interconnect_0:msgdma_tx_mm_read_readdata -> msgdma_tx:mm_read_readdata
	wire         msgdma_tx_mm_read_waitrequest;                                       // mm_interconnect_0:msgdma_tx_mm_read_waitrequest -> msgdma_tx:mm_read_waitrequest
	wire  [26:0] msgdma_tx_mm_read_address;                                           // msgdma_tx:mm_read_address -> mm_interconnect_0:msgdma_tx_mm_read_address
	wire         msgdma_tx_mm_read_read;                                              // msgdma_tx:mm_read_read -> mm_interconnect_0:msgdma_tx_mm_read_read
	wire   [3:0] msgdma_tx_mm_read_byteenable;                                        // msgdma_tx:mm_read_byteenable -> mm_interconnect_0:msgdma_tx_mm_read_byteenable
	wire         msgdma_tx_mm_read_readdatavalid;                                     // mm_interconnect_0:msgdma_tx_mm_read_readdatavalid -> msgdma_tx:mm_read_readdatavalid
	wire         msgdma_rx_mm_write_waitrequest;                                      // mm_interconnect_0:msgdma_rx_mm_write_waitrequest -> msgdma_rx:mm_write_waitrequest
	wire  [26:0] msgdma_rx_mm_write_address;                                          // msgdma_rx:mm_write_address -> mm_interconnect_0:msgdma_rx_mm_write_address
	wire   [3:0] msgdma_rx_mm_write_byteenable;                                       // msgdma_rx:mm_write_byteenable -> mm_interconnect_0:msgdma_rx_mm_write_byteenable
	wire         msgdma_rx_mm_write_write;                                            // msgdma_rx:mm_write_write -> mm_interconnect_0:msgdma_rx_mm_write_write
	wire  [31:0] msgdma_rx_mm_write_writedata;                                        // msgdma_rx:mm_write_writedata -> mm_interconnect_0:msgdma_rx_mm_write_writedata
	wire  [31:0] mm_interconnect_0_ext_epcq_flash_avl_csr_readdata;                   // ext_epcq_flash:avl_csr_rddata -> mm_interconnect_0:ext_epcq_flash_avl_csr_readdata
	wire         mm_interconnect_0_ext_epcq_flash_avl_csr_waitrequest;                // ext_epcq_flash:avl_csr_waitrequest -> mm_interconnect_0:ext_epcq_flash_avl_csr_waitrequest
	wire   [3:0] mm_interconnect_0_ext_epcq_flash_avl_csr_address;                    // mm_interconnect_0:ext_epcq_flash_avl_csr_address -> ext_epcq_flash:avl_csr_addr
	wire         mm_interconnect_0_ext_epcq_flash_avl_csr_read;                       // mm_interconnect_0:ext_epcq_flash_avl_csr_read -> ext_epcq_flash:avl_csr_read
	wire         mm_interconnect_0_ext_epcq_flash_avl_csr_readdatavalid;              // ext_epcq_flash:avl_csr_rddata_valid -> mm_interconnect_0:ext_epcq_flash_avl_csr_readdatavalid
	wire         mm_interconnect_0_ext_epcq_flash_avl_csr_write;                      // mm_interconnect_0:ext_epcq_flash_avl_csr_write -> ext_epcq_flash:avl_csr_write
	wire  [31:0] mm_interconnect_0_ext_epcq_flash_avl_csr_writedata;                  // mm_interconnect_0:ext_epcq_flash_avl_csr_writedata -> ext_epcq_flash:avl_csr_wrdata
	wire  [31:0] mm_interconnect_0_remote_update_avl_csr_readdata;                    // remote_update:avl_csr_readdata -> mm_interconnect_0:remote_update_avl_csr_readdata
	wire         mm_interconnect_0_remote_update_avl_csr_waitrequest;                 // remote_update:avl_csr_waitrequest -> mm_interconnect_0:remote_update_avl_csr_waitrequest
	wire   [4:0] mm_interconnect_0_remote_update_avl_csr_address;                     // mm_interconnect_0:remote_update_avl_csr_address -> remote_update:avl_csr_address
	wire         mm_interconnect_0_remote_update_avl_csr_read;                        // mm_interconnect_0:remote_update_avl_csr_read -> remote_update:avl_csr_read
	wire         mm_interconnect_0_remote_update_avl_csr_readdatavalid;               // remote_update:avl_csr_readdatavalid -> mm_interconnect_0:remote_update_avl_csr_readdatavalid
	wire         mm_interconnect_0_remote_update_avl_csr_write;                       // mm_interconnect_0:remote_update_avl_csr_write -> remote_update:avl_csr_write
	wire  [31:0] mm_interconnect_0_remote_update_avl_csr_writedata;                   // mm_interconnect_0:remote_update_avl_csr_writedata -> remote_update:avl_csr_writedata
	wire  [31:0] mm_interconnect_0_ext_epcq_flash_avl_mem_readdata;                   // ext_epcq_flash:avl_mem_rddata -> mm_interconnect_0:ext_epcq_flash_avl_mem_readdata
	wire         mm_interconnect_0_ext_epcq_flash_avl_mem_waitrequest;                // ext_epcq_flash:avl_mem_waitrequest -> mm_interconnect_0:ext_epcq_flash_avl_mem_waitrequest
	wire  [20:0] mm_interconnect_0_ext_epcq_flash_avl_mem_address;                    // mm_interconnect_0:ext_epcq_flash_avl_mem_address -> ext_epcq_flash:avl_mem_addr
	wire         mm_interconnect_0_ext_epcq_flash_avl_mem_read;                       // mm_interconnect_0:ext_epcq_flash_avl_mem_read -> ext_epcq_flash:avl_mem_read
	wire   [3:0] mm_interconnect_0_ext_epcq_flash_avl_mem_byteenable;                 // mm_interconnect_0:ext_epcq_flash_avl_mem_byteenable -> ext_epcq_flash:avl_mem_byteenable
	wire         mm_interconnect_0_ext_epcq_flash_avl_mem_readdatavalid;              // ext_epcq_flash:avl_mem_rddata_valid -> mm_interconnect_0:ext_epcq_flash_avl_mem_readdatavalid
	wire         mm_interconnect_0_ext_epcq_flash_avl_mem_write;                      // mm_interconnect_0:ext_epcq_flash_avl_mem_write -> ext_epcq_flash:avl_mem_write
	wire  [31:0] mm_interconnect_0_ext_epcq_flash_avl_mem_writedata;                  // mm_interconnect_0:ext_epcq_flash_avl_mem_writedata -> ext_epcq_flash:avl_mem_wrdata
	wire   [6:0] mm_interconnect_0_ext_epcq_flash_avl_mem_burstcount;                 // mm_interconnect_0:ext_epcq_flash_avl_mem_burstcount -> ext_epcq_flash:avl_mem_burstcount
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;                      // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;                   // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;                   // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;                       // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                          // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;                    // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;                         // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;                     // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_readdata;      // sll_hyperbus_controller_top_0:o_iavs0_rdata -> mm_interconnect_0:sll_hyperbus_controller_top_0_iavs0_readdata
	wire         mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_waitrequest;   // sll_hyperbus_controller_top_0:o_iavs0_wait_request -> mm_interconnect_0:sll_hyperbus_controller_top_0_iavs0_waitrequest
	wire  [21:0] mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_address;       // mm_interconnect_0:sll_hyperbus_controller_top_0_iavs0_address -> sll_hyperbus_controller_top_0:i_iavs0_addr
	wire         mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_read;          // mm_interconnect_0:sll_hyperbus_controller_top_0_iavs0_read -> sll_hyperbus_controller_top_0:i_iavs0_do_rd
	wire   [3:0] mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_byteenable;    // mm_interconnect_0:sll_hyperbus_controller_top_0_iavs0_byteenable -> sll_hyperbus_controller_top_0:i_iavs0_byteenable
	wire         mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_readdatavalid; // sll_hyperbus_controller_top_0:o_iavs0_rdata_valid -> mm_interconnect_0:sll_hyperbus_controller_top_0_iavs0_readdatavalid
	wire         mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_write;         // mm_interconnect_0:sll_hyperbus_controller_top_0_iavs0_write -> sll_hyperbus_controller_top_0:i_iavs0_do_wr
	wire  [31:0] mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_writedata;     // mm_interconnect_0:sll_hyperbus_controller_top_0_iavs0_writedata -> sll_hyperbus_controller_top_0:i_iavs0_wdata
	wire   [3:0] mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_burstcount;    // mm_interconnect_0:sll_hyperbus_controller_top_0_iavs0_burstcount -> sll_hyperbus_controller_top_0:i_iavs0_burstcount
	wire  [31:0] mm_interconnect_0_mm_bridge_0_s0_readdata;                           // mm_bridge_0:s0_readdata -> mm_interconnect_0:mm_bridge_0_s0_readdata
	wire         mm_interconnect_0_mm_bridge_0_s0_waitrequest;                        // mm_bridge_0:s0_waitrequest -> mm_interconnect_0:mm_bridge_0_s0_waitrequest
	wire         mm_interconnect_0_mm_bridge_0_s0_debugaccess;                        // mm_interconnect_0:mm_bridge_0_s0_debugaccess -> mm_bridge_0:s0_debugaccess
	wire  [14:0] mm_interconnect_0_mm_bridge_0_s0_address;                            // mm_interconnect_0:mm_bridge_0_s0_address -> mm_bridge_0:s0_address
	wire         mm_interconnect_0_mm_bridge_0_s0_read;                               // mm_interconnect_0:mm_bridge_0_s0_read -> mm_bridge_0:s0_read
	wire   [3:0] mm_interconnect_0_mm_bridge_0_s0_byteenable;                         // mm_interconnect_0:mm_bridge_0_s0_byteenable -> mm_bridge_0:s0_byteenable
	wire         mm_interconnect_0_mm_bridge_0_s0_readdatavalid;                      // mm_bridge_0:s0_readdatavalid -> mm_interconnect_0:mm_bridge_0_s0_readdatavalid
	wire         mm_interconnect_0_mm_bridge_0_s0_write;                              // mm_interconnect_0:mm_bridge_0_s0_write -> mm_bridge_0:s0_write
	wire  [31:0] mm_interconnect_0_mm_bridge_0_s0_writedata;                          // mm_interconnect_0:mm_bridge_0_s0_writedata -> mm_bridge_0:s0_writedata
	wire   [0:0] mm_interconnect_0_mm_bridge_0_s0_burstcount;                         // mm_interconnect_0:mm_bridge_0_s0_burstcount -> mm_bridge_0:s0_burstcount
	wire         mm_interconnect_0_onchip_ram_s1_chipselect;                          // mm_interconnect_0:onchip_ram_s1_chipselect -> onchip_ram:chipselect
	wire  [31:0] mm_interconnect_0_onchip_ram_s1_readdata;                            // onchip_ram:readdata -> mm_interconnect_0:onchip_ram_s1_readdata
	wire   [8:0] mm_interconnect_0_onchip_ram_s1_address;                             // mm_interconnect_0:onchip_ram_s1_address -> onchip_ram:address
	wire   [3:0] mm_interconnect_0_onchip_ram_s1_byteenable;                          // mm_interconnect_0:onchip_ram_s1_byteenable -> onchip_ram:byteenable
	wire         mm_interconnect_0_onchip_ram_s1_write;                               // mm_interconnect_0:onchip_ram_s1_write -> onchip_ram:write
	wire  [31:0] mm_interconnect_0_onchip_ram_s1_writedata;                           // mm_interconnect_0:onchip_ram_s1_writedata -> onchip_ram:writedata
	wire         mm_interconnect_0_onchip_ram_s1_clken;                               // mm_interconnect_0:onchip_ram_s1_clken -> onchip_ram:clken
	wire  [31:0] msgdma_rx_descriptor_read_master_readdata;                           // mm_interconnect_1:msgdma_rx_descriptor_read_master_readdata -> msgdma_rx:descriptor_read_master_readdata
	wire         msgdma_rx_descriptor_read_master_waitrequest;                        // mm_interconnect_1:msgdma_rx_descriptor_read_master_waitrequest -> msgdma_rx:descriptor_read_master_waitrequest
	wire  [14:0] msgdma_rx_descriptor_read_master_address;                            // msgdma_rx:descriptor_read_master_address -> mm_interconnect_1:msgdma_rx_descriptor_read_master_address
	wire         msgdma_rx_descriptor_read_master_read;                               // msgdma_rx:descriptor_read_master_read -> mm_interconnect_1:msgdma_rx_descriptor_read_master_read
	wire         msgdma_rx_descriptor_read_master_readdatavalid;                      // mm_interconnect_1:msgdma_rx_descriptor_read_master_readdatavalid -> msgdma_rx:descriptor_read_master_readdatavalid
	wire  [31:0] msgdma_tx_descriptor_read_master_readdata;                           // mm_interconnect_1:msgdma_tx_descriptor_read_master_readdata -> msgdma_tx:descriptor_read_master_readdata
	wire         msgdma_tx_descriptor_read_master_waitrequest;                        // mm_interconnect_1:msgdma_tx_descriptor_read_master_waitrequest -> msgdma_tx:descriptor_read_master_waitrequest
	wire  [14:0] msgdma_tx_descriptor_read_master_address;                            // msgdma_tx:descriptor_read_master_address -> mm_interconnect_1:msgdma_tx_descriptor_read_master_address
	wire         msgdma_tx_descriptor_read_master_read;                               // msgdma_tx:descriptor_read_master_read -> mm_interconnect_1:msgdma_tx_descriptor_read_master_read
	wire         msgdma_tx_descriptor_read_master_readdatavalid;                      // mm_interconnect_1:msgdma_tx_descriptor_read_master_readdatavalid -> msgdma_tx:descriptor_read_master_readdatavalid
	wire         msgdma_rx_descriptor_write_master_waitrequest;                       // mm_interconnect_1:msgdma_rx_descriptor_write_master_waitrequest -> msgdma_rx:descriptor_write_master_waitrequest
	wire  [14:0] msgdma_rx_descriptor_write_master_address;                           // msgdma_rx:descriptor_write_master_address -> mm_interconnect_1:msgdma_rx_descriptor_write_master_address
	wire   [3:0] msgdma_rx_descriptor_write_master_byteenable;                        // msgdma_rx:descriptor_write_master_byteenable -> mm_interconnect_1:msgdma_rx_descriptor_write_master_byteenable
	wire   [1:0] msgdma_rx_descriptor_write_master_response;                          // mm_interconnect_1:msgdma_rx_descriptor_write_master_response -> msgdma_rx:descriptor_write_master_response
	wire         msgdma_rx_descriptor_write_master_write;                             // msgdma_rx:descriptor_write_master_write -> mm_interconnect_1:msgdma_rx_descriptor_write_master_write
	wire  [31:0] msgdma_rx_descriptor_write_master_writedata;                         // msgdma_rx:descriptor_write_master_writedata -> mm_interconnect_1:msgdma_rx_descriptor_write_master_writedata
	wire         msgdma_rx_descriptor_write_master_writeresponsevalid;                // mm_interconnect_1:msgdma_rx_descriptor_write_master_writeresponsevalid -> msgdma_rx:descriptor_write_master_writeresponsevalid
	wire         msgdma_tx_descriptor_write_master_waitrequest;                       // mm_interconnect_1:msgdma_tx_descriptor_write_master_waitrequest -> msgdma_tx:descriptor_write_master_waitrequest
	wire  [14:0] msgdma_tx_descriptor_write_master_address;                           // msgdma_tx:descriptor_write_master_address -> mm_interconnect_1:msgdma_tx_descriptor_write_master_address
	wire   [3:0] msgdma_tx_descriptor_write_master_byteenable;                        // msgdma_tx:descriptor_write_master_byteenable -> mm_interconnect_1:msgdma_tx_descriptor_write_master_byteenable
	wire   [1:0] msgdma_tx_descriptor_write_master_response;                          // mm_interconnect_1:msgdma_tx_descriptor_write_master_response -> msgdma_tx:descriptor_write_master_response
	wire         msgdma_tx_descriptor_write_master_write;                             // msgdma_tx:descriptor_write_master_write -> mm_interconnect_1:msgdma_tx_descriptor_write_master_write
	wire  [31:0] msgdma_tx_descriptor_write_master_writedata;                         // msgdma_tx:descriptor_write_master_writedata -> mm_interconnect_1:msgdma_tx_descriptor_write_master_writedata
	wire         msgdma_tx_descriptor_write_master_writeresponsevalid;                // mm_interconnect_1:msgdma_tx_descriptor_write_master_writeresponsevalid -> msgdma_tx:descriptor_write_master_writeresponsevalid
	wire         mm_bridge_0_m0_waitrequest;                                          // mm_interconnect_1:mm_bridge_0_m0_waitrequest -> mm_bridge_0:m0_waitrequest
	wire  [31:0] mm_bridge_0_m0_readdata;                                             // mm_interconnect_1:mm_bridge_0_m0_readdata -> mm_bridge_0:m0_readdata
	wire         mm_bridge_0_m0_debugaccess;                                          // mm_bridge_0:m0_debugaccess -> mm_interconnect_1:mm_bridge_0_m0_debugaccess
	wire  [14:0] mm_bridge_0_m0_address;                                              // mm_bridge_0:m0_address -> mm_interconnect_1:mm_bridge_0_m0_address
	wire         mm_bridge_0_m0_read;                                                 // mm_bridge_0:m0_read -> mm_interconnect_1:mm_bridge_0_m0_read
	wire   [3:0] mm_bridge_0_m0_byteenable;                                           // mm_bridge_0:m0_byteenable -> mm_interconnect_1:mm_bridge_0_m0_byteenable
	wire         mm_bridge_0_m0_readdatavalid;                                        // mm_interconnect_1:mm_bridge_0_m0_readdatavalid -> mm_bridge_0:m0_readdatavalid
	wire  [31:0] mm_bridge_0_m0_writedata;                                            // mm_bridge_0:m0_writedata -> mm_interconnect_1:mm_bridge_0_m0_writedata
	wire         mm_bridge_0_m0_write;                                                // mm_bridge_0:m0_write -> mm_interconnect_1:mm_bridge_0_m0_write
	wire   [0:0] mm_bridge_0_m0_burstcount;                                           // mm_bridge_0:m0_burstcount -> mm_interconnect_1:mm_bridge_0_m0_burstcount
	wire         mm_interconnect_1_descriptor_memory_s1_chipselect;                   // mm_interconnect_1:descriptor_memory_s1_chipselect -> descriptor_memory:chipselect
	wire  [31:0] mm_interconnect_1_descriptor_memory_s1_readdata;                     // descriptor_memory:readdata -> mm_interconnect_1:descriptor_memory_s1_readdata
	wire  [10:0] mm_interconnect_1_descriptor_memory_s1_address;                      // mm_interconnect_1:descriptor_memory_s1_address -> descriptor_memory:address
	wire   [3:0] mm_interconnect_1_descriptor_memory_s1_byteenable;                   // mm_interconnect_1:descriptor_memory_s1_byteenable -> descriptor_memory:byteenable
	wire         mm_interconnect_1_descriptor_memory_s1_write;                        // mm_interconnect_1:descriptor_memory_s1_write -> descriptor_memory:write
	wire  [31:0] mm_interconnect_1_descriptor_memory_s1_writedata;                    // mm_interconnect_1:descriptor_memory_s1_writedata -> descriptor_memory:writedata
	wire         mm_interconnect_1_descriptor_memory_s1_clken;                        // mm_interconnect_1:descriptor_memory_s1_clken -> descriptor_memory:clken
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect;            // mm_interconnect_1:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata;              // jtag_uart:av_readdata -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest;           // jtag_uart:av_waitrequest -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_address;               // mm_interconnect_1:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_read;                  // mm_interconnect_1:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_write;                 // mm_interconnect_1:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata;             // mm_interconnect_1:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire         mm_interconnect_1_opencores_i2c_0_avalon_slave_0_chipselect;         // mm_interconnect_1:opencores_i2c_0_avalon_slave_0_chipselect -> opencores_i2c_0:wb_stb_i
	wire   [7:0] mm_interconnect_1_opencores_i2c_0_avalon_slave_0_readdata;           // opencores_i2c_0:wb_dat_o -> mm_interconnect_1:opencores_i2c_0_avalon_slave_0_readdata
	wire         mm_interconnect_1_opencores_i2c_0_avalon_slave_0_waitrequest;        // opencores_i2c_0:wb_ack_o -> mm_interconnect_1:opencores_i2c_0_avalon_slave_0_waitrequest
	wire   [2:0] mm_interconnect_1_opencores_i2c_0_avalon_slave_0_address;            // mm_interconnect_1:opencores_i2c_0_avalon_slave_0_address -> opencores_i2c_0:wb_adr_i
	wire         mm_interconnect_1_opencores_i2c_0_avalon_slave_0_write;              // mm_interconnect_1:opencores_i2c_0_avalon_slave_0_write -> opencores_i2c_0:wb_we_i
	wire   [7:0] mm_interconnect_1_opencores_i2c_0_avalon_slave_0_writedata;          // mm_interconnect_1:opencores_i2c_0_avalon_slave_0_writedata -> opencores_i2c_0:wb_dat_i
	wire  [31:0] mm_interconnect_1_eth_tse_control_port_readdata;                     // eth_tse:reg_data_out -> mm_interconnect_1:eth_tse_control_port_readdata
	wire         mm_interconnect_1_eth_tse_control_port_waitrequest;                  // eth_tse:reg_busy -> mm_interconnect_1:eth_tse_control_port_waitrequest
	wire   [7:0] mm_interconnect_1_eth_tse_control_port_address;                      // mm_interconnect_1:eth_tse_control_port_address -> eth_tse:reg_addr
	wire         mm_interconnect_1_eth_tse_control_port_read;                         // mm_interconnect_1:eth_tse_control_port_read -> eth_tse:reg_rd
	wire         mm_interconnect_1_eth_tse_control_port_write;                        // mm_interconnect_1:eth_tse_control_port_write -> eth_tse:reg_wr
	wire  [31:0] mm_interconnect_1_eth_tse_control_port_writedata;                    // mm_interconnect_1:eth_tse_control_port_writedata -> eth_tse:reg_data_in
	wire  [31:0] mm_interconnect_1_sysid_control_slave_readdata;                      // sysid:readdata -> mm_interconnect_1:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_1_sysid_control_slave_address;                       // mm_interconnect_1:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_1_msgdma_rx_csr_readdata;                            // msgdma_rx:csr_readdata -> mm_interconnect_1:msgdma_rx_csr_readdata
	wire   [2:0] mm_interconnect_1_msgdma_rx_csr_address;                             // mm_interconnect_1:msgdma_rx_csr_address -> msgdma_rx:csr_address
	wire         mm_interconnect_1_msgdma_rx_csr_read;                                // mm_interconnect_1:msgdma_rx_csr_read -> msgdma_rx:csr_read
	wire   [3:0] mm_interconnect_1_msgdma_rx_csr_byteenable;                          // mm_interconnect_1:msgdma_rx_csr_byteenable -> msgdma_rx:csr_byteenable
	wire         mm_interconnect_1_msgdma_rx_csr_write;                               // mm_interconnect_1:msgdma_rx_csr_write -> msgdma_rx:csr_write
	wire  [31:0] mm_interconnect_1_msgdma_rx_csr_writedata;                           // mm_interconnect_1:msgdma_rx_csr_writedata -> msgdma_rx:csr_writedata
	wire  [31:0] mm_interconnect_1_msgdma_tx_csr_readdata;                            // msgdma_tx:csr_readdata -> mm_interconnect_1:msgdma_tx_csr_readdata
	wire   [2:0] mm_interconnect_1_msgdma_tx_csr_address;                             // mm_interconnect_1:msgdma_tx_csr_address -> msgdma_tx:csr_address
	wire         mm_interconnect_1_msgdma_tx_csr_read;                                // mm_interconnect_1:msgdma_tx_csr_read -> msgdma_tx:csr_read
	wire   [3:0] mm_interconnect_1_msgdma_tx_csr_byteenable;                          // mm_interconnect_1:msgdma_tx_csr_byteenable -> msgdma_tx:csr_byteenable
	wire         mm_interconnect_1_msgdma_tx_csr_write;                               // mm_interconnect_1:msgdma_tx_csr_write -> msgdma_tx:csr_write
	wire  [31:0] mm_interconnect_1_msgdma_tx_csr_writedata;                           // mm_interconnect_1:msgdma_tx_csr_writedata -> msgdma_tx:csr_writedata
	wire  [31:0] mm_interconnect_1_msgdma_tx_prefetcher_csr_readdata;                 // msgdma_tx:prefetcher_csr_readdata -> mm_interconnect_1:msgdma_tx_prefetcher_csr_readdata
	wire   [2:0] mm_interconnect_1_msgdma_tx_prefetcher_csr_address;                  // mm_interconnect_1:msgdma_tx_prefetcher_csr_address -> msgdma_tx:prefetcher_csr_address
	wire         mm_interconnect_1_msgdma_tx_prefetcher_csr_read;                     // mm_interconnect_1:msgdma_tx_prefetcher_csr_read -> msgdma_tx:prefetcher_csr_read
	wire         mm_interconnect_1_msgdma_tx_prefetcher_csr_write;                    // mm_interconnect_1:msgdma_tx_prefetcher_csr_write -> msgdma_tx:prefetcher_csr_write
	wire  [31:0] mm_interconnect_1_msgdma_tx_prefetcher_csr_writedata;                // mm_interconnect_1:msgdma_tx_prefetcher_csr_writedata -> msgdma_tx:prefetcher_csr_writedata
	wire  [31:0] mm_interconnect_1_msgdma_rx_prefetcher_csr_readdata;                 // msgdma_rx:prefetcher_csr_readdata -> mm_interconnect_1:msgdma_rx_prefetcher_csr_readdata
	wire   [2:0] mm_interconnect_1_msgdma_rx_prefetcher_csr_address;                  // mm_interconnect_1:msgdma_rx_prefetcher_csr_address -> msgdma_rx:prefetcher_csr_address
	wire         mm_interconnect_1_msgdma_rx_prefetcher_csr_read;                     // mm_interconnect_1:msgdma_rx_prefetcher_csr_read -> msgdma_rx:prefetcher_csr_read
	wire         mm_interconnect_1_msgdma_rx_prefetcher_csr_write;                    // mm_interconnect_1:msgdma_rx_prefetcher_csr_write -> msgdma_rx:prefetcher_csr_write
	wire  [31:0] mm_interconnect_1_msgdma_rx_prefetcher_csr_writedata;                // mm_interconnect_1:msgdma_rx_prefetcher_csr_writedata -> msgdma_rx:prefetcher_csr_writedata
	wire         mm_interconnect_1_sys_clk_timer_s1_chipselect;                       // mm_interconnect_1:sys_clk_timer_s1_chipselect -> sys_clk_timer:chipselect
	wire  [15:0] mm_interconnect_1_sys_clk_timer_s1_readdata;                         // sys_clk_timer:readdata -> mm_interconnect_1:sys_clk_timer_s1_readdata
	wire   [2:0] mm_interconnect_1_sys_clk_timer_s1_address;                          // mm_interconnect_1:sys_clk_timer_s1_address -> sys_clk_timer:address
	wire         mm_interconnect_1_sys_clk_timer_s1_write;                            // mm_interconnect_1:sys_clk_timer_s1_write -> sys_clk_timer:write_n
	wire  [15:0] mm_interconnect_1_sys_clk_timer_s1_writedata;                        // mm_interconnect_1:sys_clk_timer_s1_writedata -> sys_clk_timer:writedata
	wire         mm_interconnect_1_led_pio_s1_chipselect;                             // mm_interconnect_1:led_pio_s1_chipselect -> led_pio:chipselect
	wire  [31:0] mm_interconnect_1_led_pio_s1_readdata;                               // led_pio:readdata -> mm_interconnect_1:led_pio_s1_readdata
	wire   [1:0] mm_interconnect_1_led_pio_s1_address;                                // mm_interconnect_1:led_pio_s1_address -> led_pio:address
	wire         mm_interconnect_1_led_pio_s1_write;                                  // mm_interconnect_1:led_pio_s1_write -> led_pio:write_n
	wire  [31:0] mm_interconnect_1_led_pio_s1_writedata;                              // mm_interconnect_1:led_pio_s1_writedata -> led_pio:writedata
	wire  [31:0] mm_interconnect_1_user_dipsw_s1_readdata;                            // user_dipsw:readdata -> mm_interconnect_1:user_dipsw_s1_readdata
	wire   [1:0] mm_interconnect_1_user_dipsw_s1_address;                             // mm_interconnect_1:user_dipsw_s1_address -> user_dipsw:address
	wire  [31:0] mm_interconnect_1_user_pb_s1_readdata;                               // user_pb:readdata -> mm_interconnect_1:user_pb_s1_readdata
	wire   [1:0] mm_interconnect_1_user_pb_s1_address;                                // mm_interconnect_1:user_pb_s1_address -> user_pb:address
	wire         irq_mapper_receiver0_irq;                                            // msgdma_rx:csr_irq_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                            // msgdma_tx:csr_irq_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                            // jtag_uart:av_irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                            // sys_clk_timer:irq -> irq_mapper:receiver3_irq
	wire  [31:0] cpu_irq_irq;                                                         // irq_mapper:sender_irq -> cpu:irq
	wire         eth_tse_receive_valid;                                               // eth_tse:ff_rx_dval -> avalon_st_adapter:in_0_valid
	wire  [31:0] eth_tse_receive_data;                                                // eth_tse:ff_rx_data -> avalon_st_adapter:in_0_data
	wire         eth_tse_receive_ready;                                               // avalon_st_adapter:in_0_ready -> eth_tse:ff_rx_rdy
	wire         eth_tse_receive_startofpacket;                                       // eth_tse:ff_rx_sop -> avalon_st_adapter:in_0_startofpacket
	wire         eth_tse_receive_endofpacket;                                         // eth_tse:ff_rx_eop -> avalon_st_adapter:in_0_endofpacket
	wire   [5:0] eth_tse_receive_error;                                               // eth_tse:rx_err -> avalon_st_adapter:in_0_error
	wire   [1:0] eth_tse_receive_empty;                                               // eth_tse:ff_rx_mod -> avalon_st_adapter:in_0_empty
	wire         avalon_st_adapter_out_0_valid;                                       // avalon_st_adapter:out_0_valid -> msgdma_rx:st_sink_valid
	wire  [31:0] avalon_st_adapter_out_0_data;                                        // avalon_st_adapter:out_0_data -> msgdma_rx:st_sink_data
	wire         avalon_st_adapter_out_0_ready;                                       // msgdma_rx:st_sink_ready -> avalon_st_adapter:out_0_ready
	wire         avalon_st_adapter_out_0_startofpacket;                               // avalon_st_adapter:out_0_startofpacket -> msgdma_rx:st_sink_startofpacket
	wire         avalon_st_adapter_out_0_endofpacket;                                 // avalon_st_adapter:out_0_endofpacket -> msgdma_rx:st_sink_endofpacket
	wire   [5:0] avalon_st_adapter_out_0_error;                                       // avalon_st_adapter:out_0_error -> msgdma_rx:st_sink_error
	wire   [1:0] avalon_st_adapter_out_0_empty;                                       // avalon_st_adapter:out_0_empty -> msgdma_rx:st_sink_empty
	wire         rst_controller_reset_out_reset;                                      // rst_controller:reset_out -> [avalon_st_adapter:in_rst_0_reset, cpu:reset_n, descriptor_memory:reset, eth_tse:reset, irq_mapper:reset, jtag_uart:rst_n, led_pio:reset_n, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, mm_interconnect_1:descriptor_memory_reset1_reset_bridge_in_reset_reset, onchip_ram:reset, rst_translator:in_reset, sys_clk_timer:reset_n, sysid:reset_n]
	wire         rst_controller_reset_out_reset_req;                                  // rst_controller:reset_req -> [cpu:reset_req, descriptor_memory:reset_req, onchip_ram:reset_req, rst_translator:reset_req_in]
	wire         cpu_debug_reset_request_reset;                                       // cpu:debug_reset_request -> rst_controller:reset_in0
	wire         rst_controller_001_reset_out_reset;                                  // rst_controller_001:reset_out -> enet_pll:reset
	wire         rst_controller_002_reset_out_reset;                                  // rst_controller_002:reset_out -> [ext_epcq_flash:reset_n, mm_interconnect_0:ext_epcq_flash_reset_reset_bridge_in_reset_reset, remote_update:reset_reset]
	wire         rst_controller_003_reset_out_reset;                                  // rst_controller_003:reset_out -> sll_hyperbus_controller_top_0:i_ext_rstn

	q_sys_cpu cpu (
		.clk                                 (sll_hyperbus_controller_top_0_o_av_out_clk_clk),    //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.d_burstcount                        (cpu_data_master_burstcount),                        //                          .burstcount
		.d_readdatavalid                     (cpu_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.i_burstcount                        (cpu_instruction_master_burstcount),                 //                          .burstcount
		.i_readdatavalid                     (cpu_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	q_sys_descriptor_memory descriptor_memory (
		.clk        (sll_hyperbus_controller_top_0_o_av_out_clk_clk),    //   clk1.clk
		.address    (mm_interconnect_1_descriptor_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_1_descriptor_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_1_descriptor_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_1_descriptor_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_1_descriptor_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_1_descriptor_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_1_descriptor_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                    // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),                //       .reset_req
		.freeze     (1'b0)                                               // (terminated)
	);

	q_sys_enet_pll enet_pll (
		.clk                (enet_clk_125m_in_clk),               //       inclk_interface.clk
		.reset              (rst_controller_001_reset_out_reset), // inclk_interface_reset.reset
		.read               (),                                   //             pll_slave.read
		.write              (),                                   //                      .write
		.address            (),                                   //                      .address
		.readdata           (),                                   //                      .readdata
		.writedata          (),                                   //                      .writedata
		.c0                 (enet_pll_c0_125m_clk),               //                    c0.clk
		.c1                 (enet_pll_c1_25m_clk),                //                    c1.clk
		.c2                 (enet_pll_c2_2m5_clk),                //                    c2.clk
		.c3                 (enet_pll_c3_125m_shift_clk),         //                    c3.clk
		.c4                 (enet_pll_c4_25m_shift_clk),          //                    c4.clk
		.areset             (enet_pll_areset_conduit_export),     //        areset_conduit.export
		.locked             (enet_pll_locked_conduit_export),     //        locked_conduit.export
		.scandone           (),                                   //           (terminated)
		.scandataout        (),                                   //           (terminated)
		.phasedone          (),                                   //           (terminated)
		.phasecounterselect (4'b0000),                            //           (terminated)
		.phaseupdown        (1'b0),                               //           (terminated)
		.phasestep          (1'b0),                               //           (terminated)
		.scanclk            (1'b0),                               //           (terminated)
		.scanclkena         (1'b0),                               //           (terminated)
		.scandata           (1'b0),                               //           (terminated)
		.configupdate       (1'b0)                                //           (terminated)
	);

	q_sys_eth_tse eth_tse (
		.clk           (sll_hyperbus_controller_top_0_o_av_out_clk_clk),     // control_port_clock_connection.clk
		.reset         (rst_controller_reset_out_reset),                     //              reset_connection.reset
		.reg_addr      (mm_interconnect_1_eth_tse_control_port_address),     //                  control_port.address
		.reg_data_out  (mm_interconnect_1_eth_tse_control_port_readdata),    //                              .readdata
		.reg_rd        (mm_interconnect_1_eth_tse_control_port_read),        //                              .read
		.reg_data_in   (mm_interconnect_1_eth_tse_control_port_writedata),   //                              .writedata
		.reg_wr        (mm_interconnect_1_eth_tse_control_port_write),       //                              .write
		.reg_busy      (mm_interconnect_1_eth_tse_control_port_waitrequest), //                              .waitrequest
		.tx_clk        (eth_tse_pcs_mac_tx_clock_connection_clk),            //   pcs_mac_tx_clock_connection.clk
		.rx_clk        (eth_tse_pcs_mac_rx_clock_connection_clk),            //   pcs_mac_rx_clock_connection.clk
		.set_10        (eth_tse_mac_status_connection_set_10),               //         mac_status_connection.set_10
		.set_1000      (eth_tse_mac_status_connection_set_1000),             //                              .set_1000
		.eth_mode      (eth_tse_mac_status_connection_eth_mode),             //                              .eth_mode
		.ena_10        (eth_tse_mac_status_connection_ena_10),               //                              .ena_10
		.rgmii_in      (eth_tse_mac_rgmii_connection_rgmii_in),              //          mac_rgmii_connection.rgmii_in
		.rgmii_out     (eth_tse_mac_rgmii_connection_rgmii_out),             //                              .rgmii_out
		.rx_control    (eth_tse_mac_rgmii_connection_rx_control),            //                              .rx_control
		.tx_control    (eth_tse_mac_rgmii_connection_tx_control),            //                              .tx_control
		.ff_rx_clk     (sll_hyperbus_controller_top_0_o_av_out_clk_clk),     //      receive_clock_connection.clk
		.ff_tx_clk     (sll_hyperbus_controller_top_0_o_av_out_clk_clk),     //     transmit_clock_connection.clk
		.ff_rx_data    (eth_tse_receive_data),                               //                       receive.data
		.ff_rx_eop     (eth_tse_receive_endofpacket),                        //                              .endofpacket
		.rx_err        (eth_tse_receive_error),                              //                              .error
		.ff_rx_mod     (eth_tse_receive_empty),                              //                              .empty
		.ff_rx_rdy     (eth_tse_receive_ready),                              //                              .ready
		.ff_rx_sop     (eth_tse_receive_startofpacket),                      //                              .startofpacket
		.ff_rx_dval    (eth_tse_receive_valid),                              //                              .valid
		.ff_tx_data    (msgdma_tx_st_source_data),                           //                      transmit.data
		.ff_tx_eop     (msgdma_tx_st_source_endofpacket),                    //                              .endofpacket
		.ff_tx_err     (msgdma_tx_st_source_error),                          //                              .error
		.ff_tx_mod     (msgdma_tx_st_source_empty),                          //                              .empty
		.ff_tx_rdy     (msgdma_tx_st_source_ready),                          //                              .ready
		.ff_tx_sop     (msgdma_tx_st_source_startofpacket),                  //                              .startofpacket
		.ff_tx_wren    (msgdma_tx_st_source_valid),                          //                              .valid
		.mdc           (eth_tse_mac_mdio_connection_mdc),                    //           mac_mdio_connection.mdc
		.mdio_in       (eth_tse_mac_mdio_connection_mdio_in),                //                              .mdio_in
		.mdio_out      (eth_tse_mac_mdio_connection_mdio_out),               //                              .mdio_out
		.mdio_oen      (eth_tse_mac_mdio_connection_mdio_oen),               //                              .mdio_oen
		.magic_wakeup  (),                                                   //           mac_misc_connection.magic_wakeup
		.magic_sleep_n (),                                                   //                              .magic_sleep_n
		.ff_tx_crc_fwd (),                                                   //                              .ff_tx_crc_fwd
		.ff_tx_septy   (),                                                   //                              .ff_tx_septy
		.tx_ff_uflow   (),                                                   //                              .tx_ff_uflow
		.ff_tx_a_full  (),                                                   //                              .ff_tx_a_full
		.ff_tx_a_empty (),                                                   //                              .ff_tx_a_empty
		.rx_err_stat   (),                                                   //                              .rx_err_stat
		.rx_frm_type   (),                                                   //                              .rx_frm_type
		.ff_rx_dsav    (),                                                   //                              .ff_rx_dsav
		.ff_rx_a_full  (),                                                   //                              .ff_rx_a_full
		.ff_rx_a_empty ()                                                    //                              .ff_rx_a_empty
	);

	q_sys_ext_epcq_flash #(
		.DEVICE_FAMILY     ("Cyclone 10 LP"),
		.ASI_WIDTH         (1),
		.CS_WIDTH          (1),
		.ADDR_WIDTH        (21),
		.ASMI_ADDR_WIDTH   (24),
		.ENABLE_4BYTE_ADDR (0),
		.CHIP_SELS         (1)
	) ext_epcq_flash (
		.avl_csr_read         (mm_interconnect_0_ext_epcq_flash_avl_csr_read),          //          avl_csr.read
		.avl_csr_waitrequest  (mm_interconnect_0_ext_epcq_flash_avl_csr_waitrequest),   //                 .waitrequest
		.avl_csr_write        (mm_interconnect_0_ext_epcq_flash_avl_csr_write),         //                 .write
		.avl_csr_addr         (mm_interconnect_0_ext_epcq_flash_avl_csr_address),       //                 .address
		.avl_csr_wrdata       (mm_interconnect_0_ext_epcq_flash_avl_csr_writedata),     //                 .writedata
		.avl_csr_rddata       (mm_interconnect_0_ext_epcq_flash_avl_csr_readdata),      //                 .readdata
		.avl_csr_rddata_valid (mm_interconnect_0_ext_epcq_flash_avl_csr_readdatavalid), //                 .readdatavalid
		.avl_mem_write        (mm_interconnect_0_ext_epcq_flash_avl_mem_write),         //          avl_mem.write
		.avl_mem_burstcount   (mm_interconnect_0_ext_epcq_flash_avl_mem_burstcount),    //                 .burstcount
		.avl_mem_waitrequest  (mm_interconnect_0_ext_epcq_flash_avl_mem_waitrequest),   //                 .waitrequest
		.avl_mem_read         (mm_interconnect_0_ext_epcq_flash_avl_mem_read),          //                 .read
		.avl_mem_addr         (mm_interconnect_0_ext_epcq_flash_avl_mem_address),       //                 .address
		.avl_mem_wrdata       (mm_interconnect_0_ext_epcq_flash_avl_mem_writedata),     //                 .writedata
		.avl_mem_rddata       (mm_interconnect_0_ext_epcq_flash_avl_mem_readdata),      //                 .readdata
		.avl_mem_rddata_valid (mm_interconnect_0_ext_epcq_flash_avl_mem_readdatavalid), //                 .readdatavalid
		.avl_mem_byteenable   (mm_interconnect_0_ext_epcq_flash_avl_mem_byteenable),    //                 .byteenable
		.irq                  (),                                                       // interrupt_sender.irq
		.clk                  (clock_bridge_0_in_clk_clk),                              //       clock_sink.clk
		.reset_n              (~rst_controller_002_reset_out_reset)                     //            reset.reset_n
	);

	q_sys_jtag_uart jtag_uart (
		.clk            (sll_hyperbus_controller_top_0_o_av_out_clk_clk),            //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver2_irq)                                   //               irq.irq
	);

	q_sys_led_pio led_pio (
		.clk        (sll_hyperbus_controller_top_0_o_av_out_clk_clk), //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_1_led_pio_s1_address),           //                  s1.address
		.write_n    (~mm_interconnect_1_led_pio_s1_write),            //                    .write_n
		.writedata  (mm_interconnect_1_led_pio_s1_writedata),         //                    .writedata
		.chipselect (mm_interconnect_1_led_pio_s1_chipselect),        //                    .chipselect
		.readdata   (mm_interconnect_1_led_pio_s1_readdata),          //                    .readdata
		.out_port   (led_pio_external_connection_export)              // external_connection.export
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (15),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_0 (
		.clk              (sll_hyperbus_controller_top_0_o_av_out_clk_clk),     //   clk.clk
		.reset            (~sll_hyperbus_controller_top_0_o_av_out_rstn_reset), // reset.reset
		.s0_waitrequest   (mm_interconnect_0_mm_bridge_0_s0_waitrequest),       //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_mm_bridge_0_s0_readdata),          //      .readdata
		.s0_readdatavalid (mm_interconnect_0_mm_bridge_0_s0_readdatavalid),     //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_mm_bridge_0_s0_burstcount),        //      .burstcount
		.s0_writedata     (mm_interconnect_0_mm_bridge_0_s0_writedata),         //      .writedata
		.s0_address       (mm_interconnect_0_mm_bridge_0_s0_address),           //      .address
		.s0_write         (mm_interconnect_0_mm_bridge_0_s0_write),             //      .write
		.s0_read          (mm_interconnect_0_mm_bridge_0_s0_read),              //      .read
		.s0_byteenable    (mm_interconnect_0_mm_bridge_0_s0_byteenable),        //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_mm_bridge_0_s0_debugaccess),       //      .debugaccess
		.m0_waitrequest   (mm_bridge_0_m0_waitrequest),                         //    m0.waitrequest
		.m0_readdata      (mm_bridge_0_m0_readdata),                            //      .readdata
		.m0_readdatavalid (mm_bridge_0_m0_readdatavalid),                       //      .readdatavalid
		.m0_burstcount    (mm_bridge_0_m0_burstcount),                          //      .burstcount
		.m0_writedata     (mm_bridge_0_m0_writedata),                           //      .writedata
		.m0_address       (mm_bridge_0_m0_address),                             //      .address
		.m0_write         (mm_bridge_0_m0_write),                               //      .write
		.m0_read          (mm_bridge_0_m0_read),                                //      .read
		.m0_byteenable    (mm_bridge_0_m0_byteenable),                          //      .byteenable
		.m0_debugaccess   (mm_bridge_0_m0_debugaccess),                         //      .debugaccess
		.s0_response      (),                                                   // (terminated)
		.m0_response      (2'b00)                                               // (terminated)
	);

	q_sys_msgdma_rx msgdma_rx (
		.mm_write_address                           (msgdma_rx_mm_write_address),                           //                mm_write.address
		.mm_write_write                             (msgdma_rx_mm_write_write),                             //                        .write
		.mm_write_byteenable                        (msgdma_rx_mm_write_byteenable),                        //                        .byteenable
		.mm_write_writedata                         (msgdma_rx_mm_write_writedata),                         //                        .writedata
		.mm_write_waitrequest                       (msgdma_rx_mm_write_waitrequest),                       //                        .waitrequest
		.descriptor_read_master_address             (msgdma_rx_descriptor_read_master_address),             //  descriptor_read_master.address
		.descriptor_read_master_read                (msgdma_rx_descriptor_read_master_read),                //                        .read
		.descriptor_read_master_readdata            (msgdma_rx_descriptor_read_master_readdata),            //                        .readdata
		.descriptor_read_master_waitrequest         (msgdma_rx_descriptor_read_master_waitrequest),         //                        .waitrequest
		.descriptor_read_master_readdatavalid       (msgdma_rx_descriptor_read_master_readdatavalid),       //                        .readdatavalid
		.descriptor_write_master_address            (msgdma_rx_descriptor_write_master_address),            // descriptor_write_master.address
		.descriptor_write_master_write              (msgdma_rx_descriptor_write_master_write),              //                        .write
		.descriptor_write_master_byteenable         (msgdma_rx_descriptor_write_master_byteenable),         //                        .byteenable
		.descriptor_write_master_writedata          (msgdma_rx_descriptor_write_master_writedata),          //                        .writedata
		.descriptor_write_master_waitrequest        (msgdma_rx_descriptor_write_master_waitrequest),        //                        .waitrequest
		.descriptor_write_master_response           (msgdma_rx_descriptor_write_master_response),           //                        .response
		.descriptor_write_master_writeresponsevalid (msgdma_rx_descriptor_write_master_writeresponsevalid), //                        .writeresponsevalid
		.clock_clk                                  (sll_hyperbus_controller_top_0_o_av_out_clk_clk),       //                   clock.clk
		.reset_n_reset_n                            (sll_hyperbus_controller_top_0_o_av_out_rstn_reset),    //                 reset_n.reset_n
		.csr_writedata                              (mm_interconnect_1_msgdma_rx_csr_writedata),            //                     csr.writedata
		.csr_write                                  (mm_interconnect_1_msgdma_rx_csr_write),                //                        .write
		.csr_byteenable                             (mm_interconnect_1_msgdma_rx_csr_byteenable),           //                        .byteenable
		.csr_readdata                               (mm_interconnect_1_msgdma_rx_csr_readdata),             //                        .readdata
		.csr_read                                   (mm_interconnect_1_msgdma_rx_csr_read),                 //                        .read
		.csr_address                                (mm_interconnect_1_msgdma_rx_csr_address),              //                        .address
		.prefetcher_csr_address                     (mm_interconnect_1_msgdma_rx_prefetcher_csr_address),   //          prefetcher_csr.address
		.prefetcher_csr_read                        (mm_interconnect_1_msgdma_rx_prefetcher_csr_read),      //                        .read
		.prefetcher_csr_write                       (mm_interconnect_1_msgdma_rx_prefetcher_csr_write),     //                        .write
		.prefetcher_csr_writedata                   (mm_interconnect_1_msgdma_rx_prefetcher_csr_writedata), //                        .writedata
		.prefetcher_csr_readdata                    (mm_interconnect_1_msgdma_rx_prefetcher_csr_readdata),  //                        .readdata
		.csr_irq_irq                                (irq_mapper_receiver0_irq),                             //                 csr_irq.irq
		.st_sink_data                               (avalon_st_adapter_out_0_data),                         //                 st_sink.data
		.st_sink_valid                              (avalon_st_adapter_out_0_valid),                        //                        .valid
		.st_sink_ready                              (avalon_st_adapter_out_0_ready),                        //                        .ready
		.st_sink_startofpacket                      (avalon_st_adapter_out_0_startofpacket),                //                        .startofpacket
		.st_sink_endofpacket                        (avalon_st_adapter_out_0_endofpacket),                  //                        .endofpacket
		.st_sink_empty                              (avalon_st_adapter_out_0_empty),                        //                        .empty
		.st_sink_error                              (avalon_st_adapter_out_0_error)                         //                        .error
	);

	q_sys_msgdma_tx msgdma_tx (
		.mm_read_address                            (msgdma_tx_mm_read_address),                            //                 mm_read.address
		.mm_read_read                               (msgdma_tx_mm_read_read),                               //                        .read
		.mm_read_byteenable                         (msgdma_tx_mm_read_byteenable),                         //                        .byteenable
		.mm_read_readdata                           (msgdma_tx_mm_read_readdata),                           //                        .readdata
		.mm_read_waitrequest                        (msgdma_tx_mm_read_waitrequest),                        //                        .waitrequest
		.mm_read_readdatavalid                      (msgdma_tx_mm_read_readdatavalid),                      //                        .readdatavalid
		.descriptor_read_master_address             (msgdma_tx_descriptor_read_master_address),             //  descriptor_read_master.address
		.descriptor_read_master_read                (msgdma_tx_descriptor_read_master_read),                //                        .read
		.descriptor_read_master_readdata            (msgdma_tx_descriptor_read_master_readdata),            //                        .readdata
		.descriptor_read_master_waitrequest         (msgdma_tx_descriptor_read_master_waitrequest),         //                        .waitrequest
		.descriptor_read_master_readdatavalid       (msgdma_tx_descriptor_read_master_readdatavalid),       //                        .readdatavalid
		.descriptor_write_master_address            (msgdma_tx_descriptor_write_master_address),            // descriptor_write_master.address
		.descriptor_write_master_write              (msgdma_tx_descriptor_write_master_write),              //                        .write
		.descriptor_write_master_byteenable         (msgdma_tx_descriptor_write_master_byteenable),         //                        .byteenable
		.descriptor_write_master_writedata          (msgdma_tx_descriptor_write_master_writedata),          //                        .writedata
		.descriptor_write_master_waitrequest        (msgdma_tx_descriptor_write_master_waitrequest),        //                        .waitrequest
		.descriptor_write_master_response           (msgdma_tx_descriptor_write_master_response),           //                        .response
		.descriptor_write_master_writeresponsevalid (msgdma_tx_descriptor_write_master_writeresponsevalid), //                        .writeresponsevalid
		.clock_clk                                  (sll_hyperbus_controller_top_0_o_av_out_clk_clk),       //                   clock.clk
		.reset_n_reset_n                            (sll_hyperbus_controller_top_0_o_av_out_rstn_reset),    //                 reset_n.reset_n
		.csr_writedata                              (mm_interconnect_1_msgdma_tx_csr_writedata),            //                     csr.writedata
		.csr_write                                  (mm_interconnect_1_msgdma_tx_csr_write),                //                        .write
		.csr_byteenable                             (mm_interconnect_1_msgdma_tx_csr_byteenable),           //                        .byteenable
		.csr_readdata                               (mm_interconnect_1_msgdma_tx_csr_readdata),             //                        .readdata
		.csr_read                                   (mm_interconnect_1_msgdma_tx_csr_read),                 //                        .read
		.csr_address                                (mm_interconnect_1_msgdma_tx_csr_address),              //                        .address
		.prefetcher_csr_address                     (mm_interconnect_1_msgdma_tx_prefetcher_csr_address),   //          prefetcher_csr.address
		.prefetcher_csr_read                        (mm_interconnect_1_msgdma_tx_prefetcher_csr_read),      //                        .read
		.prefetcher_csr_write                       (mm_interconnect_1_msgdma_tx_prefetcher_csr_write),     //                        .write
		.prefetcher_csr_writedata                   (mm_interconnect_1_msgdma_tx_prefetcher_csr_writedata), //                        .writedata
		.prefetcher_csr_readdata                    (mm_interconnect_1_msgdma_tx_prefetcher_csr_readdata),  //                        .readdata
		.csr_irq_irq                                (irq_mapper_receiver1_irq),                             //                 csr_irq.irq
		.st_source_data                             (msgdma_tx_st_source_data),                             //               st_source.data
		.st_source_valid                            (msgdma_tx_st_source_valid),                            //                        .valid
		.st_source_ready                            (msgdma_tx_st_source_ready),                            //                        .ready
		.st_source_startofpacket                    (msgdma_tx_st_source_startofpacket),                    //                        .startofpacket
		.st_source_endofpacket                      (msgdma_tx_st_source_endofpacket),                      //                        .endofpacket
		.st_source_empty                            (msgdma_tx_st_source_empty),                            //                        .empty
		.st_source_error                            (msgdma_tx_st_source_error)                             //                        .error
	);

	q_sys_onchip_ram onchip_ram (
		.clk        (sll_hyperbus_controller_top_0_o_av_out_clk_clk), //   clk1.clk
		.address    (mm_interconnect_0_onchip_ram_s1_address),        //     s1.address
		.clken      (mm_interconnect_0_onchip_ram_s1_clken),          //       .clken
		.chipselect (mm_interconnect_0_onchip_ram_s1_chipselect),     //       .chipselect
		.write      (mm_interconnect_0_onchip_ram_s1_write),          //       .write
		.readdata   (mm_interconnect_0_onchip_ram_s1_readdata),       //       .readdata
		.writedata  (mm_interconnect_0_onchip_ram_s1_writedata),      //       .writedata
		.byteenable (mm_interconnect_0_onchip_ram_s1_byteenable),     //       .byteenable
		.reset      (rst_controller_reset_out_reset),                 // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),             //       .reset_req
		.freeze     (1'b0)                                            // (terminated)
	);

	opencores_i2c #(
		.FIXED_PRESCALE (5)
	) opencores_i2c_0 (
		.wb_clk_i   (sll_hyperbus_controller_top_0_o_av_out_clk_clk),               //            clock.clk
		.wb_rst_i   (~sll_hyperbus_controller_top_0_o_av_out_rstn_reset),           //      clock_reset.reset
		.scl_pad_io (opencores_i2c_scl_pad_io),                                     //         export_0.export
		.sda_pad_io (opencores_i2c_sda_pad_io),                                     //                 .export
		.wb_adr_i   (mm_interconnect_1_opencores_i2c_0_avalon_slave_0_address),     //   avalon_slave_0.address
		.wb_dat_i   (mm_interconnect_1_opencores_i2c_0_avalon_slave_0_writedata),   //                 .writedata
		.wb_dat_o   (mm_interconnect_1_opencores_i2c_0_avalon_slave_0_readdata),    //                 .readdata
		.wb_we_i    (mm_interconnect_1_opencores_i2c_0_avalon_slave_0_write),       //                 .write
		.wb_stb_i   (mm_interconnect_1_opencores_i2c_0_avalon_slave_0_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_1_opencores_i2c_0_avalon_slave_0_waitrequest), //                 .waitrequest_n
		.wb_inta_o  ()                                                              // interrupt_sender.irq
	);

	q_sys_remote_update remote_update (
		.avl_csr_write         (mm_interconnect_0_remote_update_avl_csr_write),         // avl_csr.write
		.avl_csr_read          (mm_interconnect_0_remote_update_avl_csr_read),          //        .read
		.avl_csr_writedata     (mm_interconnect_0_remote_update_avl_csr_writedata),     //        .writedata
		.avl_csr_readdata      (mm_interconnect_0_remote_update_avl_csr_readdata),      //        .readdata
		.avl_csr_readdatavalid (mm_interconnect_0_remote_update_avl_csr_readdatavalid), //        .readdatavalid
		.avl_csr_waitrequest   (mm_interconnect_0_remote_update_avl_csr_waitrequest),   //        .waitrequest
		.avl_csr_address       (mm_interconnect_0_remote_update_avl_csr_address),       //        .address
		.clock_clk             (clock_bridge_0_in_clk_clk),                             //   clock.clk
		.reset_reset           (rst_controller_002_reset_out_reset)                     //   reset.reset
	);

	sll_hyperbus_controller_top #(
		.g_iavs0_addr_width         (22),
		.g_iavs0_data_width         (32),
		.g_iavs0_av_numsymbols      (4),
		.g_iavs0_burstcount_width   (4),
		.g_iavs0_linewrap_burst     (1),
		.g_iavs0_register_rdata     (0),
		.g_iavs0_register_wdata     (0),
		.g_include_reg_avalon       (0),
		.g_include_internal_pll     (1),
		.g_input_clk_freq_in_mhz    (50),
		.g_hyperbus_freq_in_mhz     (150),
		.g_iavs_freq_in_mhz         (75),
		.g_same_iavs_hyperbus_clk   (0),
		.g_config_rd_buffer_as_sram (1),
		.g_config_wr_buffer_as_sram (1),
		.g_device_family            ("Cyclone 10 LP"),
		.g_num_chipselect           (2),
		.g_dev0_config              (32'b00000000000000000000000000000000),
		.g_dev1_config              (32'b10001111000111110000000001000001),
		.g_dev0_timing              (32'b00000000000000000000000000000000),
		.g_dev1_timing              (32'b00000000000001100111000100100001),
		.g_include_dual_rwds_pin    (0),
		.g_dqin_rdata_width         (8)
	) sll_hyperbus_controller_top_0 (
		.in_clk               (hbus_clk_clk),                                                        //        in_clk.clk
		.i_ext_rstn           (~rst_controller_003_reset_out_reset),                                 //    i_ext_rstn.reset_n
		.i_iavs0_clk          (sll_hyperbus_controller_top_0_o_av_out_clk_clk),                      //   i_iavs0_clk.clk
		.i_iavs0_rstn         (sll_hyperbus_controller_top_0_o_av_out_rstn_reset),                   //  i_iavs0_rstn.reset_n
		.i_iavs0_addr         (mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_address),       //         iavs0.address
		.i_iavs0_burstcount   (mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_burstcount),    //              .burstcount
		.o_iavs0_wait_request (mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_waitrequest),   //              .waitrequest
		.i_iavs0_do_wr        (mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_write),         //              .write
		.i_iavs0_byteenable   (mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_byteenable),    //              .byteenable
		.i_iavs0_wdata        (mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_writedata),     //              .writedata
		.i_iavs0_do_rd        (mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_read),          //              .read
		.o_iavs0_rdata        (mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_readdata),      //              .readdata
		.o_iavs0_rdata_valid  (mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_readdatavalid), //              .readdatavalid
		.HB_RSTn              (hyperbus_controller_top_HB_RSTn),                                     //    Conduit_IO.HB_RSTn
		.HB_CLK0              (hyperbus_controller_top_HB_CLK0),                                     //              .HB_CLK0
		.HB_CLK0n             (hyperbus_controller_top_HB_CLK0n),                                    //              .HB_CLK0n
		.HB_CLK1              (hyperbus_controller_top_HB_CLK1),                                     //              .HB_CLK1
		.HB_CLK1n             (hyperbus_controller_top_HB_CLK1n),                                    //              .HB_CLK1n
		.HB_CS0n              (hyperbus_controller_top_HB_CS0n),                                     //              .HB_CS0n
		.HB_CS1n              (hyperbus_controller_top_HB_CS1n),                                     //              .HB_CS1n
		.HB_WPn               (hyperbus_controller_top_HB_WPn),                                      //              .HB_WPn
		.HB_RWDS              (hyperbus_controller_top_HB_RWDS),                                     //              .HB_RWDS
		.HB_dq                (hyperbus_controller_top_HB_dq),                                       //              .HB_dq
		.HB_RSTOn             (hyperbus_controller_top_HB_RSTOn),                                    //              .HB_RSTOn
		.HB_INTn              (hyperbus_controller_top_HB_INTn),                                     //              .HB_INTn
		.o_av_out_clk         (sll_hyperbus_controller_top_0_o_av_out_clk_clk),                      //  o_av_out_clk.clk
		.o_av_out_rstn        (sll_hyperbus_controller_top_0_o_av_out_rstn_reset),                   // o_av_out_rstn.reset_n
		.o_iavs0_resp         (),                                                                    //   (terminated)
		.i_iavsr_addr         (3'b000),                                                              //   (terminated)
		.i_iavsr_do_wr        (1'b0),                                                                //   (terminated)
		.i_iavsr_do_rd        (1'b0),                                                                //   (terminated)
		.i_iavsr_wdata        (32'b00000000000000000000000000000000),                                //   (terminated)
		.o_iavsr_rdata        ()                                                                     //   (terminated)
	);

	q_sys_sys_clk_timer sys_clk_timer (
		.clk        (sll_hyperbus_controller_top_0_o_av_out_clk_clk), //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                // reset.reset_n
		.address    (mm_interconnect_1_sys_clk_timer_s1_address),     //    s1.address
		.writedata  (mm_interconnect_1_sys_clk_timer_s1_writedata),   //      .writedata
		.readdata   (mm_interconnect_1_sys_clk_timer_s1_readdata),    //      .readdata
		.chipselect (mm_interconnect_1_sys_clk_timer_s1_chipselect),  //      .chipselect
		.write_n    (~mm_interconnect_1_sys_clk_timer_s1_write),      //      .write_n
		.irq        (irq_mapper_receiver3_irq)                        //   irq.irq
	);

	q_sys_sysid sysid (
		.clock    (sll_hyperbus_controller_top_0_o_av_out_clk_clk), //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_control_slave_address)   //              .address
	);

	q_sys_user_dipsw user_dipsw (
		.clk      (sll_hyperbus_controller_top_0_o_av_out_clk_clk),    //                 clk.clk
		.reset_n  (sll_hyperbus_controller_top_0_o_av_out_rstn_reset), //               reset.reset_n
		.address  (mm_interconnect_1_user_dipsw_s1_address),           //                  s1.address
		.readdata (mm_interconnect_1_user_dipsw_s1_readdata),          //                    .readdata
		.in_port  (user_dipsw_external_connection_export)              // external_connection.export
	);

	q_sys_user_dipsw user_pb (
		.clk      (sll_hyperbus_controller_top_0_o_av_out_clk_clk),    //                 clk.clk
		.reset_n  (sll_hyperbus_controller_top_0_o_av_out_rstn_reset), //               reset.reset_n
		.address  (mm_interconnect_1_user_pb_s1_address),              //                  s1.address
		.readdata (mm_interconnect_1_user_pb_s1_readdata),             //                    .readdata
		.in_port  (user_pb_external_connection_export)                 // external_connection.export
	);

	q_sys_mm_interconnect_0 mm_interconnect_0 (
		.clock_bridge_0_out_clk_clk                                             (clock_bridge_0_in_clk_clk),                                           //                                           clock_bridge_0_out_clk.clk
		.sll_hyperbus_controller_top_0_o_av_out_clk_clk                         (sll_hyperbus_controller_top_0_o_av_out_clk_clk),                      //                       sll_hyperbus_controller_top_0_o_av_out_clk.clk
		.cpu_reset_reset_bridge_in_reset_reset                                  (rst_controller_reset_out_reset),                                      //                                  cpu_reset_reset_bridge_in_reset.reset
		.ext_epcq_flash_reset_reset_bridge_in_reset_reset                       (rst_controller_002_reset_out_reset),                                  //                       ext_epcq_flash_reset_reset_bridge_in_reset.reset
		.sll_hyperbus_controller_top_0_i_iavs0_rstn_reset_bridge_in_reset_reset (~sll_hyperbus_controller_top_0_o_av_out_rstn_reset),                  // sll_hyperbus_controller_top_0_i_iavs0_rstn_reset_bridge_in_reset.reset
		.cpu_data_master_address                                                (cpu_data_master_address),                                             //                                                  cpu_data_master.address
		.cpu_data_master_waitrequest                                            (cpu_data_master_waitrequest),                                         //                                                                 .waitrequest
		.cpu_data_master_burstcount                                             (cpu_data_master_burstcount),                                          //                                                                 .burstcount
		.cpu_data_master_byteenable                                             (cpu_data_master_byteenable),                                          //                                                                 .byteenable
		.cpu_data_master_read                                                   (cpu_data_master_read),                                                //                                                                 .read
		.cpu_data_master_readdata                                               (cpu_data_master_readdata),                                            //                                                                 .readdata
		.cpu_data_master_readdatavalid                                          (cpu_data_master_readdatavalid),                                       //                                                                 .readdatavalid
		.cpu_data_master_write                                                  (cpu_data_master_write),                                               //                                                                 .write
		.cpu_data_master_writedata                                              (cpu_data_master_writedata),                                           //                                                                 .writedata
		.cpu_data_master_debugaccess                                            (cpu_data_master_debugaccess),                                         //                                                                 .debugaccess
		.cpu_instruction_master_address                                         (cpu_instruction_master_address),                                      //                                           cpu_instruction_master.address
		.cpu_instruction_master_waitrequest                                     (cpu_instruction_master_waitrequest),                                  //                                                                 .waitrequest
		.cpu_instruction_master_burstcount                                      (cpu_instruction_master_burstcount),                                   //                                                                 .burstcount
		.cpu_instruction_master_read                                            (cpu_instruction_master_read),                                         //                                                                 .read
		.cpu_instruction_master_readdata                                        (cpu_instruction_master_readdata),                                     //                                                                 .readdata
		.cpu_instruction_master_readdatavalid                                   (cpu_instruction_master_readdatavalid),                                //                                                                 .readdatavalid
		.msgdma_rx_mm_write_address                                             (msgdma_rx_mm_write_address),                                          //                                               msgdma_rx_mm_write.address
		.msgdma_rx_mm_write_waitrequest                                         (msgdma_rx_mm_write_waitrequest),                                      //                                                                 .waitrequest
		.msgdma_rx_mm_write_byteenable                                          (msgdma_rx_mm_write_byteenable),                                       //                                                                 .byteenable
		.msgdma_rx_mm_write_write                                               (msgdma_rx_mm_write_write),                                            //                                                                 .write
		.msgdma_rx_mm_write_writedata                                           (msgdma_rx_mm_write_writedata),                                        //                                                                 .writedata
		.msgdma_tx_mm_read_address                                              (msgdma_tx_mm_read_address),                                           //                                                msgdma_tx_mm_read.address
		.msgdma_tx_mm_read_waitrequest                                          (msgdma_tx_mm_read_waitrequest),                                       //                                                                 .waitrequest
		.msgdma_tx_mm_read_byteenable                                           (msgdma_tx_mm_read_byteenable),                                        //                                                                 .byteenable
		.msgdma_tx_mm_read_read                                                 (msgdma_tx_mm_read_read),                                              //                                                                 .read
		.msgdma_tx_mm_read_readdata                                             (msgdma_tx_mm_read_readdata),                                          //                                                                 .readdata
		.msgdma_tx_mm_read_readdatavalid                                        (msgdma_tx_mm_read_readdatavalid),                                     //                                                                 .readdatavalid
		.cpu_debug_mem_slave_address                                            (mm_interconnect_0_cpu_debug_mem_slave_address),                       //                                              cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write                                              (mm_interconnect_0_cpu_debug_mem_slave_write),                         //                                                                 .write
		.cpu_debug_mem_slave_read                                               (mm_interconnect_0_cpu_debug_mem_slave_read),                          //                                                                 .read
		.cpu_debug_mem_slave_readdata                                           (mm_interconnect_0_cpu_debug_mem_slave_readdata),                      //                                                                 .readdata
		.cpu_debug_mem_slave_writedata                                          (mm_interconnect_0_cpu_debug_mem_slave_writedata),                     //                                                                 .writedata
		.cpu_debug_mem_slave_byteenable                                         (mm_interconnect_0_cpu_debug_mem_slave_byteenable),                    //                                                                 .byteenable
		.cpu_debug_mem_slave_waitrequest                                        (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),                   //                                                                 .waitrequest
		.cpu_debug_mem_slave_debugaccess                                        (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),                   //                                                                 .debugaccess
		.ext_epcq_flash_avl_csr_address                                         (mm_interconnect_0_ext_epcq_flash_avl_csr_address),                    //                                           ext_epcq_flash_avl_csr.address
		.ext_epcq_flash_avl_csr_write                                           (mm_interconnect_0_ext_epcq_flash_avl_csr_write),                      //                                                                 .write
		.ext_epcq_flash_avl_csr_read                                            (mm_interconnect_0_ext_epcq_flash_avl_csr_read),                       //                                                                 .read
		.ext_epcq_flash_avl_csr_readdata                                        (mm_interconnect_0_ext_epcq_flash_avl_csr_readdata),                   //                                                                 .readdata
		.ext_epcq_flash_avl_csr_writedata                                       (mm_interconnect_0_ext_epcq_flash_avl_csr_writedata),                  //                                                                 .writedata
		.ext_epcq_flash_avl_csr_readdatavalid                                   (mm_interconnect_0_ext_epcq_flash_avl_csr_readdatavalid),              //                                                                 .readdatavalid
		.ext_epcq_flash_avl_csr_waitrequest                                     (mm_interconnect_0_ext_epcq_flash_avl_csr_waitrequest),                //                                                                 .waitrequest
		.ext_epcq_flash_avl_mem_address                                         (mm_interconnect_0_ext_epcq_flash_avl_mem_address),                    //                                           ext_epcq_flash_avl_mem.address
		.ext_epcq_flash_avl_mem_write                                           (mm_interconnect_0_ext_epcq_flash_avl_mem_write),                      //                                                                 .write
		.ext_epcq_flash_avl_mem_read                                            (mm_interconnect_0_ext_epcq_flash_avl_mem_read),                       //                                                                 .read
		.ext_epcq_flash_avl_mem_readdata                                        (mm_interconnect_0_ext_epcq_flash_avl_mem_readdata),                   //                                                                 .readdata
		.ext_epcq_flash_avl_mem_writedata                                       (mm_interconnect_0_ext_epcq_flash_avl_mem_writedata),                  //                                                                 .writedata
		.ext_epcq_flash_avl_mem_burstcount                                      (mm_interconnect_0_ext_epcq_flash_avl_mem_burstcount),                 //                                                                 .burstcount
		.ext_epcq_flash_avl_mem_byteenable                                      (mm_interconnect_0_ext_epcq_flash_avl_mem_byteenable),                 //                                                                 .byteenable
		.ext_epcq_flash_avl_mem_readdatavalid                                   (mm_interconnect_0_ext_epcq_flash_avl_mem_readdatavalid),              //                                                                 .readdatavalid
		.ext_epcq_flash_avl_mem_waitrequest                                     (mm_interconnect_0_ext_epcq_flash_avl_mem_waitrequest),                //                                                                 .waitrequest
		.mm_bridge_0_s0_address                                                 (mm_interconnect_0_mm_bridge_0_s0_address),                            //                                                   mm_bridge_0_s0.address
		.mm_bridge_0_s0_write                                                   (mm_interconnect_0_mm_bridge_0_s0_write),                              //                                                                 .write
		.mm_bridge_0_s0_read                                                    (mm_interconnect_0_mm_bridge_0_s0_read),                               //                                                                 .read
		.mm_bridge_0_s0_readdata                                                (mm_interconnect_0_mm_bridge_0_s0_readdata),                           //                                                                 .readdata
		.mm_bridge_0_s0_writedata                                               (mm_interconnect_0_mm_bridge_0_s0_writedata),                          //                                                                 .writedata
		.mm_bridge_0_s0_burstcount                                              (mm_interconnect_0_mm_bridge_0_s0_burstcount),                         //                                                                 .burstcount
		.mm_bridge_0_s0_byteenable                                              (mm_interconnect_0_mm_bridge_0_s0_byteenable),                         //                                                                 .byteenable
		.mm_bridge_0_s0_readdatavalid                                           (mm_interconnect_0_mm_bridge_0_s0_readdatavalid),                      //                                                                 .readdatavalid
		.mm_bridge_0_s0_waitrequest                                             (mm_interconnect_0_mm_bridge_0_s0_waitrequest),                        //                                                                 .waitrequest
		.mm_bridge_0_s0_debugaccess                                             (mm_interconnect_0_mm_bridge_0_s0_debugaccess),                        //                                                                 .debugaccess
		.onchip_ram_s1_address                                                  (mm_interconnect_0_onchip_ram_s1_address),                             //                                                    onchip_ram_s1.address
		.onchip_ram_s1_write                                                    (mm_interconnect_0_onchip_ram_s1_write),                               //                                                                 .write
		.onchip_ram_s1_readdata                                                 (mm_interconnect_0_onchip_ram_s1_readdata),                            //                                                                 .readdata
		.onchip_ram_s1_writedata                                                (mm_interconnect_0_onchip_ram_s1_writedata),                           //                                                                 .writedata
		.onchip_ram_s1_byteenable                                               (mm_interconnect_0_onchip_ram_s1_byteenable),                          //                                                                 .byteenable
		.onchip_ram_s1_chipselect                                               (mm_interconnect_0_onchip_ram_s1_chipselect),                          //                                                                 .chipselect
		.onchip_ram_s1_clken                                                    (mm_interconnect_0_onchip_ram_s1_clken),                               //                                                                 .clken
		.remote_update_avl_csr_address                                          (mm_interconnect_0_remote_update_avl_csr_address),                     //                                            remote_update_avl_csr.address
		.remote_update_avl_csr_write                                            (mm_interconnect_0_remote_update_avl_csr_write),                       //                                                                 .write
		.remote_update_avl_csr_read                                             (mm_interconnect_0_remote_update_avl_csr_read),                        //                                                                 .read
		.remote_update_avl_csr_readdata                                         (mm_interconnect_0_remote_update_avl_csr_readdata),                    //                                                                 .readdata
		.remote_update_avl_csr_writedata                                        (mm_interconnect_0_remote_update_avl_csr_writedata),                   //                                                                 .writedata
		.remote_update_avl_csr_readdatavalid                                    (mm_interconnect_0_remote_update_avl_csr_readdatavalid),               //                                                                 .readdatavalid
		.remote_update_avl_csr_waitrequest                                      (mm_interconnect_0_remote_update_avl_csr_waitrequest),                 //                                                                 .waitrequest
		.sll_hyperbus_controller_top_0_iavs0_address                            (mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_address),       //                              sll_hyperbus_controller_top_0_iavs0.address
		.sll_hyperbus_controller_top_0_iavs0_write                              (mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_write),         //                                                                 .write
		.sll_hyperbus_controller_top_0_iavs0_read                               (mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_read),          //                                                                 .read
		.sll_hyperbus_controller_top_0_iavs0_readdata                           (mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_readdata),      //                                                                 .readdata
		.sll_hyperbus_controller_top_0_iavs0_writedata                          (mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_writedata),     //                                                                 .writedata
		.sll_hyperbus_controller_top_0_iavs0_burstcount                         (mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_burstcount),    //                                                                 .burstcount
		.sll_hyperbus_controller_top_0_iavs0_byteenable                         (mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_byteenable),    //                                                                 .byteenable
		.sll_hyperbus_controller_top_0_iavs0_readdatavalid                      (mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_readdatavalid), //                                                                 .readdatavalid
		.sll_hyperbus_controller_top_0_iavs0_waitrequest                        (mm_interconnect_0_sll_hyperbus_controller_top_0_iavs0_waitrequest)    //                                                                 .waitrequest
	);

	q_sys_mm_interconnect_1 mm_interconnect_1 (
		.sll_hyperbus_controller_top_0_o_av_out_clk_clk       (sll_hyperbus_controller_top_0_o_av_out_clk_clk),                //     sll_hyperbus_controller_top_0_o_av_out_clk.clk
		.descriptor_memory_reset1_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                // descriptor_memory_reset1_reset_bridge_in_reset.reset
		.msgdma_rx_reset_n_reset_bridge_in_reset_reset        (~sll_hyperbus_controller_top_0_o_av_out_rstn_reset),            //        msgdma_rx_reset_n_reset_bridge_in_reset.reset
		.mm_bridge_0_m0_address                               (mm_bridge_0_m0_address),                                        //                                 mm_bridge_0_m0.address
		.mm_bridge_0_m0_waitrequest                           (mm_bridge_0_m0_waitrequest),                                    //                                               .waitrequest
		.mm_bridge_0_m0_burstcount                            (mm_bridge_0_m0_burstcount),                                     //                                               .burstcount
		.mm_bridge_0_m0_byteenable                            (mm_bridge_0_m0_byteenable),                                     //                                               .byteenable
		.mm_bridge_0_m0_read                                  (mm_bridge_0_m0_read),                                           //                                               .read
		.mm_bridge_0_m0_readdata                              (mm_bridge_0_m0_readdata),                                       //                                               .readdata
		.mm_bridge_0_m0_readdatavalid                         (mm_bridge_0_m0_readdatavalid),                                  //                                               .readdatavalid
		.mm_bridge_0_m0_write                                 (mm_bridge_0_m0_write),                                          //                                               .write
		.mm_bridge_0_m0_writedata                             (mm_bridge_0_m0_writedata),                                      //                                               .writedata
		.mm_bridge_0_m0_debugaccess                           (mm_bridge_0_m0_debugaccess),                                    //                                               .debugaccess
		.msgdma_rx_descriptor_read_master_address             (msgdma_rx_descriptor_read_master_address),                      //               msgdma_rx_descriptor_read_master.address
		.msgdma_rx_descriptor_read_master_waitrequest         (msgdma_rx_descriptor_read_master_waitrequest),                  //                                               .waitrequest
		.msgdma_rx_descriptor_read_master_read                (msgdma_rx_descriptor_read_master_read),                         //                                               .read
		.msgdma_rx_descriptor_read_master_readdata            (msgdma_rx_descriptor_read_master_readdata),                     //                                               .readdata
		.msgdma_rx_descriptor_read_master_readdatavalid       (msgdma_rx_descriptor_read_master_readdatavalid),                //                                               .readdatavalid
		.msgdma_rx_descriptor_write_master_address            (msgdma_rx_descriptor_write_master_address),                     //              msgdma_rx_descriptor_write_master.address
		.msgdma_rx_descriptor_write_master_waitrequest        (msgdma_rx_descriptor_write_master_waitrequest),                 //                                               .waitrequest
		.msgdma_rx_descriptor_write_master_byteenable         (msgdma_rx_descriptor_write_master_byteenable),                  //                                               .byteenable
		.msgdma_rx_descriptor_write_master_write              (msgdma_rx_descriptor_write_master_write),                       //                                               .write
		.msgdma_rx_descriptor_write_master_writedata          (msgdma_rx_descriptor_write_master_writedata),                   //                                               .writedata
		.msgdma_rx_descriptor_write_master_response           (msgdma_rx_descriptor_write_master_response),                    //                                               .response
		.msgdma_rx_descriptor_write_master_writeresponsevalid (msgdma_rx_descriptor_write_master_writeresponsevalid),          //                                               .writeresponsevalid
		.msgdma_tx_descriptor_read_master_address             (msgdma_tx_descriptor_read_master_address),                      //               msgdma_tx_descriptor_read_master.address
		.msgdma_tx_descriptor_read_master_waitrequest         (msgdma_tx_descriptor_read_master_waitrequest),                  //                                               .waitrequest
		.msgdma_tx_descriptor_read_master_read                (msgdma_tx_descriptor_read_master_read),                         //                                               .read
		.msgdma_tx_descriptor_read_master_readdata            (msgdma_tx_descriptor_read_master_readdata),                     //                                               .readdata
		.msgdma_tx_descriptor_read_master_readdatavalid       (msgdma_tx_descriptor_read_master_readdatavalid),                //                                               .readdatavalid
		.msgdma_tx_descriptor_write_master_address            (msgdma_tx_descriptor_write_master_address),                     //              msgdma_tx_descriptor_write_master.address
		.msgdma_tx_descriptor_write_master_waitrequest        (msgdma_tx_descriptor_write_master_waitrequest),                 //                                               .waitrequest
		.msgdma_tx_descriptor_write_master_byteenable         (msgdma_tx_descriptor_write_master_byteenable),                  //                                               .byteenable
		.msgdma_tx_descriptor_write_master_write              (msgdma_tx_descriptor_write_master_write),                       //                                               .write
		.msgdma_tx_descriptor_write_master_writedata          (msgdma_tx_descriptor_write_master_writedata),                   //                                               .writedata
		.msgdma_tx_descriptor_write_master_response           (msgdma_tx_descriptor_write_master_response),                    //                                               .response
		.msgdma_tx_descriptor_write_master_writeresponsevalid (msgdma_tx_descriptor_write_master_writeresponsevalid),          //                                               .writeresponsevalid
		.descriptor_memory_s1_address                         (mm_interconnect_1_descriptor_memory_s1_address),                //                           descriptor_memory_s1.address
		.descriptor_memory_s1_write                           (mm_interconnect_1_descriptor_memory_s1_write),                  //                                               .write
		.descriptor_memory_s1_readdata                        (mm_interconnect_1_descriptor_memory_s1_readdata),               //                                               .readdata
		.descriptor_memory_s1_writedata                       (mm_interconnect_1_descriptor_memory_s1_writedata),              //                                               .writedata
		.descriptor_memory_s1_byteenable                      (mm_interconnect_1_descriptor_memory_s1_byteenable),             //                                               .byteenable
		.descriptor_memory_s1_chipselect                      (mm_interconnect_1_descriptor_memory_s1_chipselect),             //                                               .chipselect
		.descriptor_memory_s1_clken                           (mm_interconnect_1_descriptor_memory_s1_clken),                  //                                               .clken
		.eth_tse_control_port_address                         (mm_interconnect_1_eth_tse_control_port_address),                //                           eth_tse_control_port.address
		.eth_tse_control_port_write                           (mm_interconnect_1_eth_tse_control_port_write),                  //                                               .write
		.eth_tse_control_port_read                            (mm_interconnect_1_eth_tse_control_port_read),                   //                                               .read
		.eth_tse_control_port_readdata                        (mm_interconnect_1_eth_tse_control_port_readdata),               //                                               .readdata
		.eth_tse_control_port_writedata                       (mm_interconnect_1_eth_tse_control_port_writedata),              //                                               .writedata
		.eth_tse_control_port_waitrequest                     (mm_interconnect_1_eth_tse_control_port_waitrequest),            //                                               .waitrequest
		.jtag_uart_avalon_jtag_slave_address                  (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),         //                    jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),           //                                               .write
		.jtag_uart_avalon_jtag_slave_read                     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),            //                                               .read
		.jtag_uart_avalon_jtag_slave_readdata                 (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),        //                                               .readdata
		.jtag_uart_avalon_jtag_slave_writedata                (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),       //                                               .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest              (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest),     //                                               .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect               (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),      //                                               .chipselect
		.led_pio_s1_address                                   (mm_interconnect_1_led_pio_s1_address),                          //                                     led_pio_s1.address
		.led_pio_s1_write                                     (mm_interconnect_1_led_pio_s1_write),                            //                                               .write
		.led_pio_s1_readdata                                  (mm_interconnect_1_led_pio_s1_readdata),                         //                                               .readdata
		.led_pio_s1_writedata                                 (mm_interconnect_1_led_pio_s1_writedata),                        //                                               .writedata
		.led_pio_s1_chipselect                                (mm_interconnect_1_led_pio_s1_chipselect),                       //                                               .chipselect
		.msgdma_rx_csr_address                                (mm_interconnect_1_msgdma_rx_csr_address),                       //                                  msgdma_rx_csr.address
		.msgdma_rx_csr_write                                  (mm_interconnect_1_msgdma_rx_csr_write),                         //                                               .write
		.msgdma_rx_csr_read                                   (mm_interconnect_1_msgdma_rx_csr_read),                          //                                               .read
		.msgdma_rx_csr_readdata                               (mm_interconnect_1_msgdma_rx_csr_readdata),                      //                                               .readdata
		.msgdma_rx_csr_writedata                              (mm_interconnect_1_msgdma_rx_csr_writedata),                     //                                               .writedata
		.msgdma_rx_csr_byteenable                             (mm_interconnect_1_msgdma_rx_csr_byteenable),                    //                                               .byteenable
		.msgdma_rx_prefetcher_csr_address                     (mm_interconnect_1_msgdma_rx_prefetcher_csr_address),            //                       msgdma_rx_prefetcher_csr.address
		.msgdma_rx_prefetcher_csr_write                       (mm_interconnect_1_msgdma_rx_prefetcher_csr_write),              //                                               .write
		.msgdma_rx_prefetcher_csr_read                        (mm_interconnect_1_msgdma_rx_prefetcher_csr_read),               //                                               .read
		.msgdma_rx_prefetcher_csr_readdata                    (mm_interconnect_1_msgdma_rx_prefetcher_csr_readdata),           //                                               .readdata
		.msgdma_rx_prefetcher_csr_writedata                   (mm_interconnect_1_msgdma_rx_prefetcher_csr_writedata),          //                                               .writedata
		.msgdma_tx_csr_address                                (mm_interconnect_1_msgdma_tx_csr_address),                       //                                  msgdma_tx_csr.address
		.msgdma_tx_csr_write                                  (mm_interconnect_1_msgdma_tx_csr_write),                         //                                               .write
		.msgdma_tx_csr_read                                   (mm_interconnect_1_msgdma_tx_csr_read),                          //                                               .read
		.msgdma_tx_csr_readdata                               (mm_interconnect_1_msgdma_tx_csr_readdata),                      //                                               .readdata
		.msgdma_tx_csr_writedata                              (mm_interconnect_1_msgdma_tx_csr_writedata),                     //                                               .writedata
		.msgdma_tx_csr_byteenable                             (mm_interconnect_1_msgdma_tx_csr_byteenable),                    //                                               .byteenable
		.msgdma_tx_prefetcher_csr_address                     (mm_interconnect_1_msgdma_tx_prefetcher_csr_address),            //                       msgdma_tx_prefetcher_csr.address
		.msgdma_tx_prefetcher_csr_write                       (mm_interconnect_1_msgdma_tx_prefetcher_csr_write),              //                                               .write
		.msgdma_tx_prefetcher_csr_read                        (mm_interconnect_1_msgdma_tx_prefetcher_csr_read),               //                                               .read
		.msgdma_tx_prefetcher_csr_readdata                    (mm_interconnect_1_msgdma_tx_prefetcher_csr_readdata),           //                                               .readdata
		.msgdma_tx_prefetcher_csr_writedata                   (mm_interconnect_1_msgdma_tx_prefetcher_csr_writedata),          //                                               .writedata
		.opencores_i2c_0_avalon_slave_0_address               (mm_interconnect_1_opencores_i2c_0_avalon_slave_0_address),      //                 opencores_i2c_0_avalon_slave_0.address
		.opencores_i2c_0_avalon_slave_0_write                 (mm_interconnect_1_opencores_i2c_0_avalon_slave_0_write),        //                                               .write
		.opencores_i2c_0_avalon_slave_0_readdata              (mm_interconnect_1_opencores_i2c_0_avalon_slave_0_readdata),     //                                               .readdata
		.opencores_i2c_0_avalon_slave_0_writedata             (mm_interconnect_1_opencores_i2c_0_avalon_slave_0_writedata),    //                                               .writedata
		.opencores_i2c_0_avalon_slave_0_waitrequest           (~mm_interconnect_1_opencores_i2c_0_avalon_slave_0_waitrequest), //                                               .waitrequest
		.opencores_i2c_0_avalon_slave_0_chipselect            (mm_interconnect_1_opencores_i2c_0_avalon_slave_0_chipselect),   //                                               .chipselect
		.sys_clk_timer_s1_address                             (mm_interconnect_1_sys_clk_timer_s1_address),                    //                               sys_clk_timer_s1.address
		.sys_clk_timer_s1_write                               (mm_interconnect_1_sys_clk_timer_s1_write),                      //                                               .write
		.sys_clk_timer_s1_readdata                            (mm_interconnect_1_sys_clk_timer_s1_readdata),                   //                                               .readdata
		.sys_clk_timer_s1_writedata                           (mm_interconnect_1_sys_clk_timer_s1_writedata),                  //                                               .writedata
		.sys_clk_timer_s1_chipselect                          (mm_interconnect_1_sys_clk_timer_s1_chipselect),                 //                                               .chipselect
		.sysid_control_slave_address                          (mm_interconnect_1_sysid_control_slave_address),                 //                            sysid_control_slave.address
		.sysid_control_slave_readdata                         (mm_interconnect_1_sysid_control_slave_readdata),                //                                               .readdata
		.user_dipsw_s1_address                                (mm_interconnect_1_user_dipsw_s1_address),                       //                                  user_dipsw_s1.address
		.user_dipsw_s1_readdata                               (mm_interconnect_1_user_dipsw_s1_readdata),                      //                                               .readdata
		.user_pb_s1_address                                   (mm_interconnect_1_user_pb_s1_address),                          //                                     user_pb_s1.address
		.user_pb_s1_readdata                                  (mm_interconnect_1_user_pb_s1_readdata)                          //                                               .readdata
	);

	q_sys_irq_mapper irq_mapper (
		.clk           (sll_hyperbus_controller_top_0_o_av_out_clk_clk), //       clk.clk
		.reset         (rst_controller_reset_out_reset),                 // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),                       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),                       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),                       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),                       // receiver3.irq
		.sender_irq    (cpu_irq_irq)                                     //    sender.irq
	);

	q_sys_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (6),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (2),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (6),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (sll_hyperbus_controller_top_0_o_av_out_clk_clk), // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),                 // in_rst_0.reset
		.in_0_data           (eth_tse_receive_data),                           //     in_0.data
		.in_0_valid          (eth_tse_receive_valid),                          //         .valid
		.in_0_ready          (eth_tse_receive_ready),                          //         .ready
		.in_0_startofpacket  (eth_tse_receive_startofpacket),                  //         .startofpacket
		.in_0_endofpacket    (eth_tse_receive_endofpacket),                    //         .endofpacket
		.in_0_empty          (eth_tse_receive_empty),                          //         .empty
		.in_0_error          (eth_tse_receive_error),                          //         .error
		.out_0_data          (avalon_st_adapter_out_0_data),                   //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),                  //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),                  //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket),          //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket),            //         .endofpacket
		.out_0_empty         (avalon_st_adapter_out_0_empty),                  //         .empty
		.out_0_error         (avalon_st_adapter_out_0_error)                   //         .error
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (cpu_debug_reset_request_reset),                      // reset_in0.reset
		.reset_in1      (~sll_hyperbus_controller_top_0_o_av_out_rstn_reset), // reset_in1.reset
		.clk            (sll_hyperbus_controller_top_0_o_av_out_clk_clk),     //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),                     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),                 //          .reset_req
		.reset_req_in0  (1'b0),                                               // (terminated)
		.reset_req_in1  (1'b0),                                               // (terminated)
		.reset_in2      (1'b0),                                               // (terminated)
		.reset_req_in2  (1'b0),                                               // (terminated)
		.reset_in3      (1'b0),                                               // (terminated)
		.reset_req_in3  (1'b0),                                               // (terminated)
		.reset_in4      (1'b0),                                               // (terminated)
		.reset_req_in4  (1'b0),                                               // (terminated)
		.reset_in5      (1'b0),                                               // (terminated)
		.reset_req_in5  (1'b0),                                               // (terminated)
		.reset_in6      (1'b0),                                               // (terminated)
		.reset_req_in6  (1'b0),                                               // (terminated)
		.reset_in7      (1'b0),                                               // (terminated)
		.reset_req_in7  (1'b0),                                               // (terminated)
		.reset_in8      (1'b0),                                               // (terminated)
		.reset_req_in8  (1'b0),                                               // (terminated)
		.reset_in9      (1'b0),                                               // (terminated)
		.reset_req_in9  (1'b0),                                               // (terminated)
		.reset_in10     (1'b0),                                               // (terminated)
		.reset_req_in10 (1'b0),                                               // (terminated)
		.reset_in11     (1'b0),                                               // (terminated)
		.reset_req_in11 (1'b0),                                               // (terminated)
		.reset_in12     (1'b0),                                               // (terminated)
		.reset_req_in12 (1'b0),                                               // (terminated)
		.reset_in13     (1'b0),                                               // (terminated)
		.reset_req_in13 (1'b0),                                               // (terminated)
		.reset_in14     (1'b0),                                               // (terminated)
		.reset_req_in14 (1'b0),                                               // (terminated)
		.reset_in15     (1'b0),                                               // (terminated)
		.reset_req_in15 (1'b0)                                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_enet_reset_n),                // reset_in0.reset
		.clk            (enet_clk_125m_in_clk),               //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~hbus_reset_reset_n),                // reset_in0.reset
		.clk            (clock_bridge_0_in_clk_clk),          //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~hbus_reset_reset_n),                // reset_in0.reset
		.clk            (hbus_clk_clk),                       //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
